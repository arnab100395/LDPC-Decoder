module Ldpc_Decoder_final(clk,reset,L1,L2,L3,L4,L5,L6,L7,L8,L9,L10,L11,L12,L13,L14,L15,L16,L17,L18,L19,L20,L21,L22,L23,L24,L25,L26,L27,L28,L29,L30,L31,L32,L33,L34,L35,L36,L37,L38,L39,L40,L41,L42,L43,L44,L45,L46,L47,L48,L49,L50,L51,L52,L53,L54,L55,L56,L57,L58,L59,L60,L61,L62,L63,L64,L65,L66,L67,L68,L69,L70,L71,L72,L73,L74,L75,L76,L77,L78,L79,L80,L81,L82,L83,L84,L85,L86,L87,L88,L89,L90,L91,L92,L93,L94,L95,L96,L97,L98,L99,L100,L101,L102,L103,L104,L105,L106,L107,L108,L109,L110,L111,L112,L113,L114,L115,L116,L117,L118,L119,L120,L121,L122,L123,L124,L125,L126,L127,L128,L129,L130,L131,L132,L133,L134,L135,L136,L137,L138,L139,L140,L141,L142,L143,L144,L145,L146,L147,L148,L149,L150,L151,L152,L153,L154,L155,L156,L157,L158,L159,L160,L161,L162,L163,L164,L165,L166,L167,L168,L169,L170,L171,L172,L173,L174,L175,L176,L177,L178,L179,L180,L181,L182,L183,L184,L185,L186,L187,L188,L189,L190,L191,L192,L193,L194,L195,L196,L197,L198,L199,L200,L201,L202,L203,L204,L205,L206,L207,L208,L209,L210,L211,L212,L213,L214,L215,L216,L217,L218,L219,L220,L221,L222,L223,L224,L225,L226,L227,L228,L229,L230,L231,L232,L233,L234,L235,L236,L237,L238,L239,L240,L241,L242,L243,L244,L245,L246,L247,L248,L249,L250,L251,L252,L253,L254,L255,L256,L257,L258,L259,L260,L261,L262,L263,L264,L265,L266,L267,L268,L269,L270,L271,L272,L273,L274,L275,L276,L277,L278,L279,L280,L281,L282,L283,L284,L285,L286,L287,L288,L289,L290,L291,L292,L293,L294,L295,L296,L297,L298,L299,L300,L301,L302,L303,L304,L305,L306,L307,L308,L309,L310,L311,L312,L313,L314,L315,L316,L317,L318,L319,L320,L321,L322,L323,L324,L325,L326,L327,L328,L329,L330,L331,L332,L333,L334,L335,L336,L337,L338,L339,L340,L341,L342,L343,L344,L345,L346,L347,L348,L349,L350,L351,L352,L353,L354,L355,L356,L357,L358,L359,L360,L361,L362,L363,L364,L365,L366,L367,L368,L369,L370,L371,L372,L373,L374,L375,L376,L377,L378,L379,L380,L381,L382,L383,L384,L385,L386,L387,L388,L389,L390,L391,L392,L393,L394,L395,L396,L397,L398,L399,L400,L401,L402,L403,L404,L405,L406,L407,L408,L409,L410,L411,L412,L413,L414,L415,L416,L417,L418,L419,L420,L421,L422,L423,L424,L425,L426,L427,L428,L429,L430,L431,L432,L433,L434,L435,L436,L437,L438,L439,L440,L441,L442,L443,L444,L445,L446,L447,L448,L449,L450,L451,L452,L453,L454,L455,L456,L457,L458,L459,L460,L461,L462,L463,L464,L465,L466,L467,L468,L469,L470,L471,L472,L473,L474,L475,L476,L477,L478,L479,L480,L481,L482,L483,L484,L485,L486,L487,L488,L489,L490,L491,L492,L493,L494,L495,L496,L497,L498,L499,L500,L501,L502,L503,L504,L505,L506,L507,L508,L509,L510,L511,L512,L513,L514,L515,L516,L517,L518,L519,L520,L521,L522,L523,L524,L525,L526,L527,L528,L529,L530,L531,L532,L533,L534,L535,L536,L537,L538,L539,L540,L541,L542,L543,L544,L545,L546,L547,L548,L549,L550,L551,L552,L553,L554,L555,L556,L557,L558,L559,L560,L561,L562,L563,L564,L565,L566,L567,L568,L569,L570,L571,L572,L573,L574,L575,L576,P);

input clk,reset;
input signed [31:0] L1,L2,L3,L4,L5,L6,L7,L8,L9,L10,L11,L12,L13,L14,L15,L16,L17,L18,L19,L20,L21,L22,L23,L24,L25,L26,L27,L28,L29,L30,L31,L32,L33,L34,L35,L36,L37,L38,L39,L40,L41,L42,L43,L44,L45,L46,L47,L48,L49,L50,L51,L52,L53,L54,L55,L56,L57,L58,L59,L60,L61,L62,L63,L64,L65,L66,L67,L68,L69,L70,L71,L72,L73,L74,L75,L76,L77,L78,L79,L80,L81,L82,L83,L84,L85,L86,L87,L88,L89,L90,L91,L92,L93,L94,L95,L96,L97,L98,L99,L100,L101,L102,L103,L104,L105,L106,L107,L108,L109,L110,L111,L112,L113,L114,L115,L116,L117,L118,L119,L120,L121,L122,L123,L124,L125,L126,L127,L128,L129,L130,L131,L132,L133,L134,L135,L136,L137,L138,L139,L140,L141,L142,L143,L144,L145,L146,L147,L148,L149,L150,L151,L152,L153,L154,L155,L156,L157,L158,L159,L160,L161,L162,L163,L164,L165,L166,L167,L168,L169,L170,L171,L172,L173,L174,L175,L176,L177,L178,L179,L180,L181,L182,L183,L184,L185,L186,L187,L188,L189,L190,L191,L192,L193,L194,L195,L196,L197,L198,L199,L200,L201,L202,L203,L204,L205,L206,L207,L208,L209,L210,L211,L212,L213,L214,L215,L216,L217,L218,L219,L220,L221,L222,L223,L224,L225,L226,L227,L228,L229,L230,L231,L232,L233,L234,L235,L236,L237,L238,L239,L240,L241,L242,L243,L244,L245,L246,L247,L248,L249,L250,L251,L252,L253,L254,L255,L256,L257,L258,L259,L260,L261,L262,L263,L264,L265,L266,L267,L268,L269,L270,L271,L272,L273,L274,L275,L276,L277,L278,L279,L280,L281,L282,L283,L284,L285,L286,L287,L288,L289,L290,L291,L292,L293,L294,L295,L296,L297,L298,L299,L300,L301,L302,L303,L304,L305,L306,L307,L308,L309,L310,L311,L312,L313,L314,L315,L316,L317,L318,L319,L320,L321,L322,L323,L324,L325,L326,L327,L328,L329,L330,L331,L332,L333,L334,L335,L336,L337,L338,L339,L340,L341,L342,L343,L344,L345,L346,L347,L348,L349,L350,L351,L352,L353,L354,L355,L356,L357,L358,L359,L360,L361,L362,L363,L364,L365,L366,L367,L368,L369,L370,L371,L372,L373,L374,L375,L376,L377,L378,L379,L380,L381,L382,L383,L384,L385,L386,L387,L388,L389,L390,L391,L392,L393,L394,L395,L396,L397,L398,L399,L400,L401,L402,L403,L404,L405,L406,L407,L408,L409,L410,L411,L412,L413,L414,L415,L416,L417,L418,L419,L420,L421,L422,L423,L424,L425,L426,L427,L428,L429,L430,L431,L432,L433,L434,L435,L436,L437,L438,L439,L440,L441,L442,L443,L444,L445,L446,L447,L448,L449,L450,L451,L452,L453,L454,L455,L456,L457,L458,L459,L460,L461,L462,L463,L464,L465,L466,L467,L468,L469,L470,L471,L472,L473,L474,L475,L476,L477,L478,L479,L480,L481,L482,L483,L484,L485,L486,L487,L488,L489,L490,L491,L492,L493,L494,L495,L496,L497,L498,L499,L500,L501,L502,L503,L504,L505,L506,L507,L508,L509,L510,L511,L512,L513,L514,L515,L516,L517,L518,L519,L520,L521,L522,L523,L524,L525,L526,L527,L528,L529,L530,L531,L532,L533,L534,L535,L536,L537,L538,L539,L540,L541,L542,L543,L544,L545,L546,L547,L548,L549,L550,L551,L552,L553,L554,L555,L556,L557,L558,L559,L560,L561,L562,L563,L564,L565,L566,L567,L568,L569,L570,L571,L572,L573,L574,L575,L576;
output [0:575] P;
wire signed [31:0] R [0:1823];
wire signed [31:0] Q [0:1823];

CNU_6 CNU1	(.Q1(Q[0])	,.Q2(Q[1])	,.Q3(Q[2])	,.Q4(Q[3])	,.Q5(Q[4])	,.Q6(Q[5])			,.R1(R[0])	,.R2(R[1])	,.R3(R[2])	,.R4(R[3])	,.R5(R[4])	,.R6(R[5])			,.clk(clk)	);
CNU_6 CNU2	(.Q1(Q[6])	,.Q2(Q[7])	,.Q3(Q[8])	,.Q4(Q[9])	,.Q5(Q[10])	,.Q6(Q[11])			,.R1(R[6])	,.R2(R[7])	,.R3(R[8])	,.R4(R[9])	,.R5(R[10])	,.R6(R[11])			,.clk(clk)	);
CNU_6 CNU3	(.Q1(Q[12])	,.Q2(Q[13])	,.Q3(Q[14])	,.Q4(Q[15])	,.Q5(Q[16])	,.Q6(Q[17])			,.R1(R[12])	,.R2(R[13])	,.R3(R[14])	,.R4(R[15])	,.R5(R[16])	,.R6(R[17])			,.clk(clk)	);
CNU_6 CNU4	(.Q1(Q[18])	,.Q2(Q[19])	,.Q3(Q[20])	,.Q4(Q[21])	,.Q5(Q[22])	,.Q6(Q[23])			,.R1(R[18])	,.R2(R[19])	,.R3(R[20])	,.R4(R[21])	,.R5(R[22])	,.R6(R[23])			,.clk(clk)	);
CNU_6 CNU5	(.Q1(Q[24])	,.Q2(Q[25])	,.Q3(Q[26])	,.Q4(Q[27])	,.Q5(Q[28])	,.Q6(Q[29])			,.R1(R[24])	,.R2(R[25])	,.R3(R[26])	,.R4(R[27])	,.R5(R[28])	,.R6(R[29])			,.clk(clk)	);
CNU_6 CNU6	(.Q1(Q[30])	,.Q2(Q[31])	,.Q3(Q[32])	,.Q4(Q[33])	,.Q5(Q[34])	,.Q6(Q[35])			,.R1(R[30])	,.R2(R[31])	,.R3(R[32])	,.R4(R[33])	,.R5(R[34])	,.R6(R[35])			,.clk(clk)	);
CNU_6 CNU7	(.Q1(Q[36])	,.Q2(Q[37])	,.Q3(Q[38])	,.Q4(Q[39])	,.Q5(Q[40])	,.Q6(Q[41])			,.R1(R[36])	,.R2(R[37])	,.R3(R[38])	,.R4(R[39])	,.R5(R[40])	,.R6(R[41])			,.clk(clk)	);
CNU_6 CNU8	(.Q1(Q[42])	,.Q2(Q[43])	,.Q3(Q[44])	,.Q4(Q[45])	,.Q5(Q[46])	,.Q6(Q[47])			,.R1(R[42])	,.R2(R[43])	,.R3(R[44])	,.R4(R[45])	,.R5(R[46])	,.R6(R[47])			,.clk(clk)	);
CNU_6 CNU9	(.Q1(Q[48])	,.Q2(Q[49])	,.Q3(Q[50])	,.Q4(Q[51])	,.Q5(Q[52])	,.Q6(Q[53])			,.R1(R[48])	,.R2(R[49])	,.R3(R[50])	,.R4(R[51])	,.R5(R[52])	,.R6(R[53])			,.clk(clk)	);
CNU_6 CNU10	(.Q1(Q[54])	,.Q2(Q[55])	,.Q3(Q[56])	,.Q4(Q[57])	,.Q5(Q[58])	,.Q6(Q[59])			,.R1(R[54])	,.R2(R[55])	,.R3(R[56])	,.R4(R[57])	,.R5(R[58])	,.R6(R[59])			,.clk(clk)	);
CNU_6 CNU11	(.Q1(Q[60])	,.Q2(Q[61])	,.Q3(Q[62])	,.Q4(Q[63])	,.Q5(Q[64])	,.Q6(Q[65])			,.R1(R[60])	,.R2(R[61])	,.R3(R[62])	,.R4(R[63])	,.R5(R[64])	,.R6(R[65])			,.clk(clk)	);
CNU_6 CNU12	(.Q1(Q[66])	,.Q2(Q[67])	,.Q3(Q[68])	,.Q4(Q[69])	,.Q5(Q[70])	,.Q6(Q[71])			,.R1(R[66])	,.R2(R[67])	,.R3(R[68])	,.R4(R[69])	,.R5(R[70])	,.R6(R[71])			,.clk(clk)	);
CNU_6 CNU13	(.Q1(Q[72])	,.Q2(Q[73])	,.Q3(Q[74])	,.Q4(Q[75])	,.Q5(Q[76])	,.Q6(Q[77])			,.R1(R[72])	,.R2(R[73])	,.R3(R[74])	,.R4(R[75])	,.R5(R[76])	,.R6(R[77])			,.clk(clk)	);
CNU_6 CNU14	(.Q1(Q[78])	,.Q2(Q[79])	,.Q3(Q[80])	,.Q4(Q[81])	,.Q5(Q[82])	,.Q6(Q[83])			,.R1(R[78])	,.R2(R[79])	,.R3(R[80])	,.R4(R[81])	,.R5(R[82])	,.R6(R[83])			,.clk(clk)	);
CNU_6 CNU15	(.Q1(Q[84])	,.Q2(Q[85])	,.Q3(Q[86])	,.Q4(Q[87])	,.Q5(Q[88])	,.Q6(Q[89])			,.R1(R[84])	,.R2(R[85])	,.R3(R[86])	,.R4(R[87])	,.R5(R[88])	,.R6(R[89])			,.clk(clk)	);
CNU_6 CNU16	(.Q1(Q[90])	,.Q2(Q[91])	,.Q3(Q[92])	,.Q4(Q[93])	,.Q5(Q[94])	,.Q6(Q[95])			,.R1(R[90])	,.R2(R[91])	,.R3(R[92])	,.R4(R[93])	,.R5(R[94])	,.R6(R[95])			,.clk(clk)	);
CNU_6 CNU17	(.Q1(Q[96])	,.Q2(Q[97])	,.Q3(Q[98])	,.Q4(Q[99])	,.Q5(Q[100])	,.Q6(Q[101])			,.R1(R[96])	,.R2(R[97])	,.R3(R[98])	,.R4(R[99])	,.R5(R[100])	,.R6(R[101])			,.clk(clk)	);
CNU_6 CNU18	(.Q1(Q[102])	,.Q2(Q[103])	,.Q3(Q[104])	,.Q4(Q[105])	,.Q5(Q[106])	,.Q6(Q[107])			,.R1(R[102])	,.R2(R[103])	,.R3(R[104])	,.R4(R[105])	,.R5(R[106])	,.R6(R[107])			,.clk(clk)	);
CNU_6 CNU19	(.Q1(Q[108])	,.Q2(Q[109])	,.Q3(Q[110])	,.Q4(Q[111])	,.Q5(Q[112])	,.Q6(Q[113])			,.R1(R[108])	,.R2(R[109])	,.R3(R[110])	,.R4(R[111])	,.R5(R[112])	,.R6(R[113])			,.clk(clk)	);
CNU_6 CNU20	(.Q1(Q[114])	,.Q2(Q[115])	,.Q3(Q[116])	,.Q4(Q[117])	,.Q5(Q[118])	,.Q6(Q[119])			,.R1(R[114])	,.R2(R[115])	,.R3(R[116])	,.R4(R[117])	,.R5(R[118])	,.R6(R[119])			,.clk(clk)	);
CNU_6 CNU21	(.Q1(Q[120])	,.Q2(Q[121])	,.Q3(Q[122])	,.Q4(Q[123])	,.Q5(Q[124])	,.Q6(Q[125])			,.R1(R[120])	,.R2(R[121])	,.R3(R[122])	,.R4(R[123])	,.R5(R[124])	,.R6(R[125])			,.clk(clk)	);
CNU_6 CNU22	(.Q1(Q[126])	,.Q2(Q[127])	,.Q3(Q[128])	,.Q4(Q[129])	,.Q5(Q[130])	,.Q6(Q[131])			,.R1(R[126])	,.R2(R[127])	,.R3(R[128])	,.R4(R[129])	,.R5(R[130])	,.R6(R[131])			,.clk(clk)	);
CNU_6 CNU23	(.Q1(Q[132])	,.Q2(Q[133])	,.Q3(Q[134])	,.Q4(Q[135])	,.Q5(Q[136])	,.Q6(Q[137])			,.R1(R[132])	,.R2(R[133])	,.R3(R[134])	,.R4(R[135])	,.R5(R[136])	,.R6(R[137])			,.clk(clk)	);
CNU_6 CNU24	(.Q1(Q[138])	,.Q2(Q[139])	,.Q3(Q[140])	,.Q4(Q[141])	,.Q5(Q[142])	,.Q6(Q[143])			,.R1(R[138])	,.R2(R[139])	,.R3(R[140])	,.R4(R[141])	,.R5(R[142])	,.R6(R[143])			,.clk(clk)	);

CNU_7 CNU25	(.Q1(Q[144])	,.Q2(Q[145])	,.Q3(Q[146])	,.Q4(Q[147])	,.Q5(Q[148])	,.Q6(Q[149])	,.Q7(Q[150])	,.R1(R[144])	,.R2(R[145])	,.R3(R[146])	,.R4(R[147])	,.R5(R[148])	,.R6(R[149])	,.R7(R[150])	,.clk(clk)	);
CNU_7 CNU26	(.Q1(Q[151])	,.Q2(Q[152])	,.Q3(Q[153])	,.Q4(Q[154])	,.Q5(Q[155])	,.Q6(Q[156])	,.Q7(Q[157])	,.R1(R[151])	,.R2(R[152])	,.R3(R[153])	,.R4(R[154])	,.R5(R[155])	,.R6(R[156])	,.R7(R[157])	,.clk(clk)	);
CNU_7 CNU27	(.Q1(Q[158])	,.Q2(Q[159])	,.Q3(Q[160])	,.Q4(Q[161])	,.Q5(Q[162])	,.Q6(Q[163])	,.Q7(Q[164])	,.R1(R[158])	,.R2(R[159])	,.R3(R[160])	,.R4(R[161])	,.R5(R[162])	,.R6(R[163])	,.R7(R[164])	,.clk(clk)	);
CNU_7 CNU28	(.Q1(Q[165])	,.Q2(Q[166])	,.Q3(Q[167])	,.Q4(Q[168])	,.Q5(Q[169])	,.Q6(Q[170])	,.Q7(Q[171])	,.R1(R[165])	,.R2(R[166])	,.R3(R[167])	,.R4(R[168])	,.R5(R[169])	,.R6(R[170])	,.R7(R[171])	,.clk(clk)	);
CNU_7 CNU29	(.Q1(Q[172])	,.Q2(Q[173])	,.Q3(Q[174])	,.Q4(Q[175])	,.Q5(Q[176])	,.Q6(Q[177])	,.Q7(Q[178])	,.R1(R[172])	,.R2(R[173])	,.R3(R[174])	,.R4(R[175])	,.R5(R[176])	,.R6(R[177])	,.R7(R[178])	,.clk(clk)	);
CNU_7 CNU30	(.Q1(Q[179])	,.Q2(Q[180])	,.Q3(Q[181])	,.Q4(Q[182])	,.Q5(Q[183])	,.Q6(Q[184])	,.Q7(Q[185])	,.R1(R[179])	,.R2(R[180])	,.R3(R[181])	,.R4(R[182])	,.R5(R[183])	,.R6(R[184])	,.R7(R[185])	,.clk(clk)	);
CNU_7 CNU31	(.Q1(Q[186])	,.Q2(Q[187])	,.Q3(Q[188])	,.Q4(Q[189])	,.Q5(Q[190])	,.Q6(Q[191])	,.Q7(Q[192])	,.R1(R[186])	,.R2(R[187])	,.R3(R[188])	,.R4(R[189])	,.R5(R[190])	,.R6(R[191])	,.R7(R[192])	,.clk(clk)	);
CNU_7 CNU32	(.Q1(Q[193])	,.Q2(Q[194])	,.Q3(Q[195])	,.Q4(Q[196])	,.Q5(Q[197])	,.Q6(Q[198])	,.Q7(Q[199])	,.R1(R[193])	,.R2(R[194])	,.R3(R[195])	,.R4(R[196])	,.R5(R[197])	,.R6(R[198])	,.R7(R[199])	,.clk(clk)	);
CNU_7 CNU33	(.Q1(Q[200])	,.Q2(Q[201])	,.Q3(Q[202])	,.Q4(Q[203])	,.Q5(Q[204])	,.Q6(Q[205])	,.Q7(Q[206])	,.R1(R[200])	,.R2(R[201])	,.R3(R[202])	,.R4(R[203])	,.R5(R[204])	,.R6(R[205])	,.R7(R[206])	,.clk(clk)	);
CNU_7 CNU34	(.Q1(Q[207])	,.Q2(Q[208])	,.Q3(Q[209])	,.Q4(Q[210])	,.Q5(Q[211])	,.Q6(Q[212])	,.Q7(Q[213])	,.R1(R[207])	,.R2(R[208])	,.R3(R[209])	,.R4(R[210])	,.R5(R[211])	,.R6(R[212])	,.R7(R[213])	,.clk(clk)	);
CNU_7 CNU35	(.Q1(Q[214])	,.Q2(Q[215])	,.Q3(Q[216])	,.Q4(Q[217])	,.Q5(Q[218])	,.Q6(Q[219])	,.Q7(Q[220])	,.R1(R[214])	,.R2(R[215])	,.R3(R[216])	,.R4(R[217])	,.R5(R[218])	,.R6(R[219])	,.R7(R[220])	,.clk(clk)	);
CNU_7 CNU36	(.Q1(Q[221])	,.Q2(Q[222])	,.Q3(Q[223])	,.Q4(Q[224])	,.Q5(Q[225])	,.Q6(Q[226])	,.Q7(Q[227])	,.R1(R[221])	,.R2(R[222])	,.R3(R[223])	,.R4(R[224])	,.R5(R[225])	,.R6(R[226])	,.R7(R[227])	,.clk(clk)	);
CNU_7 CNU37	(.Q1(Q[228])	,.Q2(Q[229])	,.Q3(Q[230])	,.Q4(Q[231])	,.Q5(Q[232])	,.Q6(Q[233])	,.Q7(Q[234])	,.R1(R[228])	,.R2(R[229])	,.R3(R[230])	,.R4(R[231])	,.R5(R[232])	,.R6(R[233])	,.R7(R[234])	,.clk(clk)	);
CNU_7 CNU38	(.Q1(Q[235])	,.Q2(Q[236])	,.Q3(Q[237])	,.Q4(Q[238])	,.Q5(Q[239])	,.Q6(Q[240])	,.Q7(Q[241])	,.R1(R[235])	,.R2(R[236])	,.R3(R[237])	,.R4(R[238])	,.R5(R[239])	,.R6(R[240])	,.R7(R[241])	,.clk(clk)	);
CNU_7 CNU39	(.Q1(Q[242])	,.Q2(Q[243])	,.Q3(Q[244])	,.Q4(Q[245])	,.Q5(Q[246])	,.Q6(Q[247])	,.Q7(Q[248])	,.R1(R[242])	,.R2(R[243])	,.R3(R[244])	,.R4(R[245])	,.R5(R[246])	,.R6(R[247])	,.R7(R[248])	,.clk(clk)	);
CNU_7 CNU40	(.Q1(Q[249])	,.Q2(Q[250])	,.Q3(Q[251])	,.Q4(Q[252])	,.Q5(Q[253])	,.Q6(Q[254])	,.Q7(Q[255])	,.R1(R[249])	,.R2(R[250])	,.R3(R[251])	,.R4(R[252])	,.R5(R[253])	,.R6(R[254])	,.R7(R[255])	,.clk(clk)	);
CNU_7 CNU41	(.Q1(Q[256])	,.Q2(Q[257])	,.Q3(Q[258])	,.Q4(Q[259])	,.Q5(Q[260])	,.Q6(Q[261])	,.Q7(Q[262])	,.R1(R[256])	,.R2(R[257])	,.R3(R[258])	,.R4(R[259])	,.R5(R[260])	,.R6(R[261])	,.R7(R[262])	,.clk(clk)	);
CNU_7 CNU42	(.Q1(Q[263])	,.Q2(Q[264])	,.Q3(Q[265])	,.Q4(Q[266])	,.Q5(Q[267])	,.Q6(Q[268])	,.Q7(Q[269])	,.R1(R[263])	,.R2(R[264])	,.R3(R[265])	,.R4(R[266])	,.R5(R[267])	,.R6(R[268])	,.R7(R[269])	,.clk(clk)	);
CNU_7 CNU43	(.Q1(Q[270])	,.Q2(Q[271])	,.Q3(Q[272])	,.Q4(Q[273])	,.Q5(Q[274])	,.Q6(Q[275])	,.Q7(Q[276])	,.R1(R[270])	,.R2(R[271])	,.R3(R[272])	,.R4(R[273])	,.R5(R[274])	,.R6(R[275])	,.R7(R[276])	,.clk(clk)	);
CNU_7 CNU44	(.Q1(Q[277])	,.Q2(Q[278])	,.Q3(Q[279])	,.Q4(Q[280])	,.Q5(Q[281])	,.Q6(Q[282])	,.Q7(Q[283])	,.R1(R[277])	,.R2(R[278])	,.R3(R[279])	,.R4(R[280])	,.R5(R[281])	,.R6(R[282])	,.R7(R[283])	,.clk(clk)	);
CNU_7 CNU45	(.Q1(Q[284])	,.Q2(Q[285])	,.Q3(Q[286])	,.Q4(Q[287])	,.Q5(Q[288])	,.Q6(Q[289])	,.Q7(Q[290])	,.R1(R[284])	,.R2(R[285])	,.R3(R[286])	,.R4(R[287])	,.R5(R[288])	,.R6(R[289])	,.R7(R[290])	,.clk(clk)	);
CNU_7 CNU46	(.Q1(Q[291])	,.Q2(Q[292])	,.Q3(Q[293])	,.Q4(Q[294])	,.Q5(Q[295])	,.Q6(Q[296])	,.Q7(Q[297])	,.R1(R[291])	,.R2(R[292])	,.R3(R[293])	,.R4(R[294])	,.R5(R[295])	,.R6(R[296])	,.R7(R[297])	,.clk(clk)	);
CNU_7 CNU47	(.Q1(Q[298])	,.Q2(Q[299])	,.Q3(Q[300])	,.Q4(Q[301])	,.Q5(Q[302])	,.Q6(Q[303])	,.Q7(Q[304])	,.R1(R[298])	,.R2(R[299])	,.R3(R[300])	,.R4(R[301])	,.R5(R[302])	,.R6(R[303])	,.R7(R[304])	,.clk(clk)	);
CNU_7 CNU48	(.Q1(Q[305])	,.Q2(Q[306])	,.Q3(Q[307])	,.Q4(Q[308])	,.Q5(Q[309])	,.Q6(Q[310])	,.Q7(Q[311])	,.R1(R[305])	,.R2(R[306])	,.R3(R[307])	,.R4(R[308])	,.R5(R[309])	,.R6(R[310])	,.R7(R[311])	,.clk(clk)	);
CNU_7 CNU49	(.Q1(Q[312])	,.Q2(Q[313])	,.Q3(Q[314])	,.Q4(Q[315])	,.Q5(Q[316])	,.Q6(Q[317])	,.Q7(Q[318])	,.R1(R[312])	,.R2(R[313])	,.R3(R[314])	,.R4(R[315])	,.R5(R[316])	,.R6(R[317])	,.R7(R[318])	,.clk(clk)	);
CNU_7 CNU50	(.Q1(Q[319])	,.Q2(Q[320])	,.Q3(Q[321])	,.Q4(Q[322])	,.Q5(Q[323])	,.Q6(Q[324])	,.Q7(Q[325])	,.R1(R[319])	,.R2(R[320])	,.R3(R[321])	,.R4(R[322])	,.R5(R[323])	,.R6(R[324])	,.R7(R[325])	,.clk(clk)	);
CNU_7 CNU51	(.Q1(Q[326])	,.Q2(Q[327])	,.Q3(Q[328])	,.Q4(Q[329])	,.Q5(Q[330])	,.Q6(Q[331])	,.Q7(Q[332])	,.R1(R[326])	,.R2(R[327])	,.R3(R[328])	,.R4(R[329])	,.R5(R[330])	,.R6(R[331])	,.R7(R[332])	,.clk(clk)	);
CNU_7 CNU52	(.Q1(Q[333])	,.Q2(Q[334])	,.Q3(Q[335])	,.Q4(Q[336])	,.Q5(Q[337])	,.Q6(Q[338])	,.Q7(Q[339])	,.R1(R[333])	,.R2(R[334])	,.R3(R[335])	,.R4(R[336])	,.R5(R[337])	,.R6(R[338])	,.R7(R[339])	,.clk(clk)	);
CNU_7 CNU53	(.Q1(Q[340])	,.Q2(Q[341])	,.Q3(Q[342])	,.Q4(Q[343])	,.Q5(Q[344])	,.Q6(Q[345])	,.Q7(Q[346])	,.R1(R[340])	,.R2(R[341])	,.R3(R[342])	,.R4(R[343])	,.R5(R[344])	,.R6(R[345])	,.R7(R[346])	,.clk(clk)	);
CNU_7 CNU54	(.Q1(Q[347])	,.Q2(Q[348])	,.Q3(Q[349])	,.Q4(Q[350])	,.Q5(Q[351])	,.Q6(Q[352])	,.Q7(Q[353])	,.R1(R[347])	,.R2(R[348])	,.R3(R[349])	,.R4(R[350])	,.R5(R[351])	,.R6(R[352])	,.R7(R[353])	,.clk(clk)	);
CNU_7 CNU55	(.Q1(Q[354])	,.Q2(Q[355])	,.Q3(Q[356])	,.Q4(Q[357])	,.Q5(Q[358])	,.Q6(Q[359])	,.Q7(Q[360])	,.R1(R[354])	,.R2(R[355])	,.R3(R[356])	,.R4(R[357])	,.R5(R[358])	,.R6(R[359])	,.R7(R[360])	,.clk(clk)	);
CNU_7 CNU56	(.Q1(Q[361])	,.Q2(Q[362])	,.Q3(Q[363])	,.Q4(Q[364])	,.Q5(Q[365])	,.Q6(Q[366])	,.Q7(Q[367])	,.R1(R[361])	,.R2(R[362])	,.R3(R[363])	,.R4(R[364])	,.R5(R[365])	,.R6(R[366])	,.R7(R[367])	,.clk(clk)	);
CNU_7 CNU57	(.Q1(Q[368])	,.Q2(Q[369])	,.Q3(Q[370])	,.Q4(Q[371])	,.Q5(Q[372])	,.Q6(Q[373])	,.Q7(Q[374])	,.R1(R[368])	,.R2(R[369])	,.R3(R[370])	,.R4(R[371])	,.R5(R[372])	,.R6(R[373])	,.R7(R[374])	,.clk(clk)	);
CNU_7 CNU58	(.Q1(Q[375])	,.Q2(Q[376])	,.Q3(Q[377])	,.Q4(Q[378])	,.Q5(Q[379])	,.Q6(Q[380])	,.Q7(Q[381])	,.R1(R[375])	,.R2(R[376])	,.R3(R[377])	,.R4(R[378])	,.R5(R[379])	,.R6(R[380])	,.R7(R[381])	,.clk(clk)	);
CNU_7 CNU59	(.Q1(Q[382])	,.Q2(Q[383])	,.Q3(Q[384])	,.Q4(Q[385])	,.Q5(Q[386])	,.Q6(Q[387])	,.Q7(Q[388])	,.R1(R[382])	,.R2(R[383])	,.R3(R[384])	,.R4(R[385])	,.R5(R[386])	,.R6(R[387])	,.R7(R[388])	,.clk(clk)	);
CNU_7 CNU60	(.Q1(Q[389])	,.Q2(Q[390])	,.Q3(Q[391])	,.Q4(Q[392])	,.Q5(Q[393])	,.Q6(Q[394])	,.Q7(Q[395])	,.R1(R[389])	,.R2(R[390])	,.R3(R[391])	,.R4(R[392])	,.R5(R[393])	,.R6(R[394])	,.R7(R[395])	,.clk(clk)	);
CNU_7 CNU61	(.Q1(Q[396])	,.Q2(Q[397])	,.Q3(Q[398])	,.Q4(Q[399])	,.Q5(Q[400])	,.Q6(Q[401])	,.Q7(Q[402])	,.R1(R[396])	,.R2(R[397])	,.R3(R[398])	,.R4(R[399])	,.R5(R[400])	,.R6(R[401])	,.R7(R[402])	,.clk(clk)	);
CNU_7 CNU62	(.Q1(Q[403])	,.Q2(Q[404])	,.Q3(Q[405])	,.Q4(Q[406])	,.Q5(Q[407])	,.Q6(Q[408])	,.Q7(Q[409])	,.R1(R[403])	,.R2(R[404])	,.R3(R[405])	,.R4(R[406])	,.R5(R[407])	,.R6(R[408])	,.R7(R[409])	,.clk(clk)	);
CNU_7 CNU63	(.Q1(Q[410])	,.Q2(Q[411])	,.Q3(Q[412])	,.Q4(Q[413])	,.Q5(Q[414])	,.Q6(Q[415])	,.Q7(Q[416])	,.R1(R[410])	,.R2(R[411])	,.R3(R[412])	,.R4(R[413])	,.R5(R[414])	,.R6(R[415])	,.R7(R[416])	,.clk(clk)	);
CNU_7 CNU64	(.Q1(Q[417])	,.Q2(Q[418])	,.Q3(Q[419])	,.Q4(Q[420])	,.Q5(Q[421])	,.Q6(Q[422])	,.Q7(Q[423])	,.R1(R[417])	,.R2(R[418])	,.R3(R[419])	,.R4(R[420])	,.R5(R[421])	,.R6(R[422])	,.R7(R[423])	,.clk(clk)	);
CNU_7 CNU65	(.Q1(Q[424])	,.Q2(Q[425])	,.Q3(Q[426])	,.Q4(Q[427])	,.Q5(Q[428])	,.Q6(Q[429])	,.Q7(Q[430])	,.R1(R[424])	,.R2(R[425])	,.R3(R[426])	,.R4(R[427])	,.R5(R[428])	,.R6(R[429])	,.R7(R[430])	,.clk(clk)	);
CNU_7 CNU66	(.Q1(Q[431])	,.Q2(Q[432])	,.Q3(Q[433])	,.Q4(Q[434])	,.Q5(Q[435])	,.Q6(Q[436])	,.Q7(Q[437])	,.R1(R[431])	,.R2(R[432])	,.R3(R[433])	,.R4(R[434])	,.R5(R[435])	,.R6(R[436])	,.R7(R[437])	,.clk(clk)	);
CNU_7 CNU67	(.Q1(Q[438])	,.Q2(Q[439])	,.Q3(Q[440])	,.Q4(Q[441])	,.Q5(Q[442])	,.Q6(Q[443])	,.Q7(Q[444])	,.R1(R[438])	,.R2(R[439])	,.R3(R[440])	,.R4(R[441])	,.R5(R[442])	,.R6(R[443])	,.R7(R[444])	,.clk(clk)	);
CNU_7 CNU68	(.Q1(Q[445])	,.Q2(Q[446])	,.Q3(Q[447])	,.Q4(Q[448])	,.Q5(Q[449])	,.Q6(Q[450])	,.Q7(Q[451])	,.R1(R[445])	,.R2(R[446])	,.R3(R[447])	,.R4(R[448])	,.R5(R[449])	,.R6(R[450])	,.R7(R[451])	,.clk(clk)	);
CNU_7 CNU69	(.Q1(Q[452])	,.Q2(Q[453])	,.Q3(Q[454])	,.Q4(Q[455])	,.Q5(Q[456])	,.Q6(Q[457])	,.Q7(Q[458])	,.R1(R[452])	,.R2(R[453])	,.R3(R[454])	,.R4(R[455])	,.R5(R[456])	,.R6(R[457])	,.R7(R[458])	,.clk(clk)	);
CNU_7 CNU70	(.Q1(Q[459])	,.Q2(Q[460])	,.Q3(Q[461])	,.Q4(Q[462])	,.Q5(Q[463])	,.Q6(Q[464])	,.Q7(Q[465])	,.R1(R[459])	,.R2(R[460])	,.R3(R[461])	,.R4(R[462])	,.R5(R[463])	,.R6(R[464])	,.R7(R[465])	,.clk(clk)	);
CNU_7 CNU71	(.Q1(Q[466])	,.Q2(Q[467])	,.Q3(Q[468])	,.Q4(Q[469])	,.Q5(Q[470])	,.Q6(Q[471])	,.Q7(Q[472])	,.R1(R[466])	,.R2(R[467])	,.R3(R[468])	,.R4(R[469])	,.R5(R[470])	,.R6(R[471])	,.R7(R[472])	,.clk(clk)	);
CNU_7 CNU72	(.Q1(Q[473])	,.Q2(Q[474])	,.Q3(Q[475])	,.Q4(Q[476])	,.Q5(Q[477])	,.Q6(Q[478])	,.Q7(Q[479])	,.R1(R[473])	,.R2(R[474])	,.R3(R[475])	,.R4(R[476])	,.R5(R[477])	,.R6(R[478])	,.R7(R[479])	,.clk(clk)	);

CNU_6 CNU73	(.Q1(Q[480])	,.Q2(Q[481])	,.Q3(Q[482])	,.Q4(Q[483])	,.Q5(Q[484])	,.Q6(Q[485])			,.R1(R[480])	,.R2(R[481])	,.R3(R[482])	,.R4(R[483])	,.R5(R[484])	,.R6(R[485])			,.clk(clk)	);
CNU_6 CNU74	(.Q1(Q[486])	,.Q2(Q[487])	,.Q3(Q[488])	,.Q4(Q[489])	,.Q5(Q[490])	,.Q6(Q[491])			,.R1(R[486])	,.R2(R[487])	,.R3(R[488])	,.R4(R[489])	,.R5(R[490])	,.R6(R[491])			,.clk(clk)	);
CNU_6 CNU75	(.Q1(Q[492])	,.Q2(Q[493])	,.Q3(Q[494])	,.Q4(Q[495])	,.Q5(Q[496])	,.Q6(Q[497])			,.R1(R[492])	,.R2(R[493])	,.R3(R[494])	,.R4(R[495])	,.R5(R[496])	,.R6(R[497])			,.clk(clk)	);
CNU_6 CNU76	(.Q1(Q[498])	,.Q2(Q[499])	,.Q3(Q[500])	,.Q4(Q[501])	,.Q5(Q[502])	,.Q6(Q[503])			,.R1(R[498])	,.R2(R[499])	,.R3(R[500])	,.R4(R[501])	,.R5(R[502])	,.R6(R[503])			,.clk(clk)	);
CNU_6 CNU77	(.Q1(Q[504])	,.Q2(Q[505])	,.Q3(Q[506])	,.Q4(Q[507])	,.Q5(Q[508])	,.Q6(Q[509])			,.R1(R[504])	,.R2(R[505])	,.R3(R[506])	,.R4(R[507])	,.R5(R[508])	,.R6(R[509])			,.clk(clk)	);
CNU_6 CNU78	(.Q1(Q[510])	,.Q2(Q[511])	,.Q3(Q[512])	,.Q4(Q[513])	,.Q5(Q[514])	,.Q6(Q[515])			,.R1(R[510])	,.R2(R[511])	,.R3(R[512])	,.R4(R[513])	,.R5(R[514])	,.R6(R[515])			,.clk(clk)	);
CNU_6 CNU79	(.Q1(Q[516])	,.Q2(Q[517])	,.Q3(Q[518])	,.Q4(Q[519])	,.Q5(Q[520])	,.Q6(Q[521])			,.R1(R[516])	,.R2(R[517])	,.R3(R[518])	,.R4(R[519])	,.R5(R[520])	,.R6(R[521])			,.clk(clk)	);
CNU_6 CNU80	(.Q1(Q[522])	,.Q2(Q[523])	,.Q3(Q[524])	,.Q4(Q[525])	,.Q5(Q[526])	,.Q6(Q[527])			,.R1(R[522])	,.R2(R[523])	,.R3(R[524])	,.R4(R[525])	,.R5(R[526])	,.R6(R[527])			,.clk(clk)	);
CNU_6 CNU81	(.Q1(Q[528])	,.Q2(Q[529])	,.Q3(Q[530])	,.Q4(Q[531])	,.Q5(Q[532])	,.Q6(Q[533])			,.R1(R[528])	,.R2(R[529])	,.R3(R[530])	,.R4(R[531])	,.R5(R[532])	,.R6(R[533])			,.clk(clk)	);
CNU_6 CNU82	(.Q1(Q[534])	,.Q2(Q[535])	,.Q3(Q[536])	,.Q4(Q[537])	,.Q5(Q[538])	,.Q6(Q[539])			,.R1(R[534])	,.R2(R[535])	,.R3(R[536])	,.R4(R[537])	,.R5(R[538])	,.R6(R[539])			,.clk(clk)	);
CNU_6 CNU83	(.Q1(Q[540])	,.Q2(Q[541])	,.Q3(Q[542])	,.Q4(Q[543])	,.Q5(Q[544])	,.Q6(Q[545])			,.R1(R[540])	,.R2(R[541])	,.R3(R[542])	,.R4(R[543])	,.R5(R[544])	,.R6(R[545])			,.clk(clk)	);
CNU_6 CNU84	(.Q1(Q[546])	,.Q2(Q[547])	,.Q3(Q[548])	,.Q4(Q[549])	,.Q5(Q[550])	,.Q6(Q[551])			,.R1(R[546])	,.R2(R[547])	,.R3(R[548])	,.R4(R[549])	,.R5(R[550])	,.R6(R[551])			,.clk(clk)	);
CNU_6 CNU85	(.Q1(Q[552])	,.Q2(Q[553])	,.Q3(Q[554])	,.Q4(Q[555])	,.Q5(Q[556])	,.Q6(Q[557])			,.R1(R[552])	,.R2(R[553])	,.R3(R[554])	,.R4(R[555])	,.R5(R[556])	,.R6(R[557])			,.clk(clk)	);
CNU_6 CNU86	(.Q1(Q[558])	,.Q2(Q[559])	,.Q3(Q[560])	,.Q4(Q[561])	,.Q5(Q[562])	,.Q6(Q[563])			,.R1(R[558])	,.R2(R[559])	,.R3(R[560])	,.R4(R[561])	,.R5(R[562])	,.R6(R[563])			,.clk(clk)	);
CNU_6 CNU87	(.Q1(Q[564])	,.Q2(Q[565])	,.Q3(Q[566])	,.Q4(Q[567])	,.Q5(Q[568])	,.Q6(Q[569])			,.R1(R[564])	,.R2(R[565])	,.R3(R[566])	,.R4(R[567])	,.R5(R[568])	,.R6(R[569])			,.clk(clk)	);
CNU_6 CNU88	(.Q1(Q[570])	,.Q2(Q[571])	,.Q3(Q[572])	,.Q4(Q[573])	,.Q5(Q[574])	,.Q6(Q[575])			,.R1(R[570])	,.R2(R[571])	,.R3(R[572])	,.R4(R[573])	,.R5(R[574])	,.R6(R[575])			,.clk(clk)	);
CNU_6 CNU89	(.Q1(Q[576])	,.Q2(Q[577])	,.Q3(Q[578])	,.Q4(Q[579])	,.Q5(Q[580])	,.Q6(Q[581])			,.R1(R[576])	,.R2(R[577])	,.R3(R[578])	,.R4(R[579])	,.R5(R[580])	,.R6(R[581])			,.clk(clk)	);
CNU_6 CNU90	(.Q1(Q[582])	,.Q2(Q[583])	,.Q3(Q[584])	,.Q4(Q[585])	,.Q5(Q[586])	,.Q6(Q[587])			,.R1(R[582])	,.R2(R[583])	,.R3(R[584])	,.R4(R[585])	,.R5(R[586])	,.R6(R[587])			,.clk(clk)	);
CNU_6 CNU91	(.Q1(Q[588])	,.Q2(Q[589])	,.Q3(Q[590])	,.Q4(Q[591])	,.Q5(Q[592])	,.Q6(Q[593])			,.R1(R[588])	,.R2(R[589])	,.R3(R[590])	,.R4(R[591])	,.R5(R[592])	,.R6(R[593])			,.clk(clk)	);
CNU_6 CNU92	(.Q1(Q[594])	,.Q2(Q[595])	,.Q3(Q[596])	,.Q4(Q[597])	,.Q5(Q[598])	,.Q6(Q[599])			,.R1(R[594])	,.R2(R[595])	,.R3(R[596])	,.R4(R[597])	,.R5(R[598])	,.R6(R[599])			,.clk(clk)	);
CNU_6 CNU93	(.Q1(Q[600])	,.Q2(Q[601])	,.Q3(Q[602])	,.Q4(Q[603])	,.Q5(Q[604])	,.Q6(Q[605])			,.R1(R[600])	,.R2(R[601])	,.R3(R[602])	,.R4(R[603])	,.R5(R[604])	,.R6(R[605])			,.clk(clk)	);
CNU_6 CNU94	(.Q1(Q[606])	,.Q2(Q[607])	,.Q3(Q[608])	,.Q4(Q[609])	,.Q5(Q[610])	,.Q6(Q[611])			,.R1(R[606])	,.R2(R[607])	,.R3(R[608])	,.R4(R[609])	,.R5(R[610])	,.R6(R[611])			,.clk(clk)	);
CNU_6 CNU95	(.Q1(Q[612])	,.Q2(Q[613])	,.Q3(Q[614])	,.Q4(Q[615])	,.Q5(Q[616])	,.Q6(Q[617])			,.R1(R[612])	,.R2(R[613])	,.R3(R[614])	,.R4(R[615])	,.R5(R[616])	,.R6(R[617])			,.clk(clk)	);
CNU_6 CNU96	(.Q1(Q[618])	,.Q2(Q[619])	,.Q3(Q[620])	,.Q4(Q[621])	,.Q5(Q[622])	,.Q6(Q[623])			,.R1(R[618])	,.R2(R[619])	,.R3(R[620])	,.R4(R[621])	,.R5(R[622])	,.R6(R[623])			,.clk(clk)	);
CNU_6 CNU97	(.Q1(Q[624])	,.Q2(Q[625])	,.Q3(Q[626])	,.Q4(Q[627])	,.Q5(Q[628])	,.Q6(Q[629])			,.R1(R[624])	,.R2(R[625])	,.R3(R[626])	,.R4(R[627])	,.R5(R[628])	,.R6(R[629])			,.clk(clk)	);
CNU_6 CNU98	(.Q1(Q[630])	,.Q2(Q[631])	,.Q3(Q[632])	,.Q4(Q[633])	,.Q5(Q[634])	,.Q6(Q[635])			,.R1(R[630])	,.R2(R[631])	,.R3(R[632])	,.R4(R[633])	,.R5(R[634])	,.R6(R[635])			,.clk(clk)	);
CNU_6 CNU99	(.Q1(Q[636])	,.Q2(Q[637])	,.Q3(Q[638])	,.Q4(Q[639])	,.Q5(Q[640])	,.Q6(Q[641])			,.R1(R[636])	,.R2(R[637])	,.R3(R[638])	,.R4(R[639])	,.R5(R[640])	,.R6(R[641])			,.clk(clk)	);
CNU_6 CNU100	(.Q1(Q[642])	,.Q2(Q[643])	,.Q3(Q[644])	,.Q4(Q[645])	,.Q5(Q[646])	,.Q6(Q[647])			,.R1(R[642])	,.R2(R[643])	,.R3(R[644])	,.R4(R[645])	,.R5(R[646])	,.R6(R[647])			,.clk(clk)	);
CNU_6 CNU101	(.Q1(Q[648])	,.Q2(Q[649])	,.Q3(Q[650])	,.Q4(Q[651])	,.Q5(Q[652])	,.Q6(Q[653])			,.R1(R[648])	,.R2(R[649])	,.R3(R[650])	,.R4(R[651])	,.R5(R[652])	,.R6(R[653])			,.clk(clk)	);
CNU_6 CNU102	(.Q1(Q[654])	,.Q2(Q[655])	,.Q3(Q[656])	,.Q4(Q[657])	,.Q5(Q[658])	,.Q6(Q[659])			,.R1(R[654])	,.R2(R[655])	,.R3(R[656])	,.R4(R[657])	,.R5(R[658])	,.R6(R[659])			,.clk(clk)	);
CNU_6 CNU103	(.Q1(Q[660])	,.Q2(Q[661])	,.Q3(Q[662])	,.Q4(Q[663])	,.Q5(Q[664])	,.Q6(Q[665])			,.R1(R[660])	,.R2(R[661])	,.R3(R[662])	,.R4(R[663])	,.R5(R[664])	,.R6(R[665])			,.clk(clk)	);
CNU_6 CNU104	(.Q1(Q[666])	,.Q2(Q[667])	,.Q3(Q[668])	,.Q4(Q[669])	,.Q5(Q[670])	,.Q6(Q[671])			,.R1(R[666])	,.R2(R[667])	,.R3(R[668])	,.R4(R[669])	,.R5(R[670])	,.R6(R[671])			,.clk(clk)	);
CNU_6 CNU105	(.Q1(Q[672])	,.Q2(Q[673])	,.Q3(Q[674])	,.Q4(Q[675])	,.Q5(Q[676])	,.Q6(Q[677])			,.R1(R[672])	,.R2(R[673])	,.R3(R[674])	,.R4(R[675])	,.R5(R[676])	,.R6(R[677])			,.clk(clk)	);
CNU_6 CNU106	(.Q1(Q[678])	,.Q2(Q[679])	,.Q3(Q[680])	,.Q4(Q[681])	,.Q5(Q[682])	,.Q6(Q[683])			,.R1(R[678])	,.R2(R[679])	,.R3(R[680])	,.R4(R[681])	,.R5(R[682])	,.R6(R[683])			,.clk(clk)	);
CNU_6 CNU107	(.Q1(Q[684])	,.Q2(Q[685])	,.Q3(Q[686])	,.Q4(Q[687])	,.Q5(Q[688])	,.Q6(Q[689])			,.R1(R[684])	,.R2(R[685])	,.R3(R[686])	,.R4(R[687])	,.R5(R[688])	,.R6(R[689])			,.clk(clk)	);
CNU_6 CNU108	(.Q1(Q[690])	,.Q2(Q[691])	,.Q3(Q[692])	,.Q4(Q[693])	,.Q5(Q[694])	,.Q6(Q[695])			,.R1(R[690])	,.R2(R[691])	,.R3(R[692])	,.R4(R[693])	,.R5(R[694])	,.R6(R[695])			,.clk(clk)	);
CNU_6 CNU109	(.Q1(Q[696])	,.Q2(Q[697])	,.Q3(Q[698])	,.Q4(Q[699])	,.Q5(Q[700])	,.Q6(Q[701])			,.R1(R[696])	,.R2(R[697])	,.R3(R[698])	,.R4(R[699])	,.R5(R[700])	,.R6(R[701])			,.clk(clk)	);
CNU_6 CNU110	(.Q1(Q[702])	,.Q2(Q[703])	,.Q3(Q[704])	,.Q4(Q[705])	,.Q5(Q[706])	,.Q6(Q[707])			,.R1(R[702])	,.R2(R[703])	,.R3(R[704])	,.R4(R[705])	,.R5(R[706])	,.R6(R[707])			,.clk(clk)	);
CNU_6 CNU111	(.Q1(Q[708])	,.Q2(Q[709])	,.Q3(Q[710])	,.Q4(Q[711])	,.Q5(Q[712])	,.Q6(Q[713])			,.R1(R[708])	,.R2(R[709])	,.R3(R[710])	,.R4(R[711])	,.R5(R[712])	,.R6(R[713])			,.clk(clk)	);
CNU_6 CNU112	(.Q1(Q[714])	,.Q2(Q[715])	,.Q3(Q[716])	,.Q4(Q[717])	,.Q5(Q[718])	,.Q6(Q[719])			,.R1(R[714])	,.R2(R[715])	,.R3(R[716])	,.R4(R[717])	,.R5(R[718])	,.R6(R[719])			,.clk(clk)	);
CNU_6 CNU113	(.Q1(Q[720])	,.Q2(Q[721])	,.Q3(Q[722])	,.Q4(Q[723])	,.Q5(Q[724])	,.Q6(Q[725])			,.R1(R[720])	,.R2(R[721])	,.R3(R[722])	,.R4(R[723])	,.R5(R[724])	,.R6(R[725])			,.clk(clk)	);
CNU_6 CNU114	(.Q1(Q[726])	,.Q2(Q[727])	,.Q3(Q[728])	,.Q4(Q[729])	,.Q5(Q[730])	,.Q6(Q[731])			,.R1(R[726])	,.R2(R[727])	,.R3(R[728])	,.R4(R[729])	,.R5(R[730])	,.R6(R[731])			,.clk(clk)	);
CNU_6 CNU115	(.Q1(Q[732])	,.Q2(Q[733])	,.Q3(Q[734])	,.Q4(Q[735])	,.Q5(Q[736])	,.Q6(Q[737])			,.R1(R[732])	,.R2(R[733])	,.R3(R[734])	,.R4(R[735])	,.R5(R[736])	,.R6(R[737])			,.clk(clk)	);
CNU_6 CNU116	(.Q1(Q[738])	,.Q2(Q[739])	,.Q3(Q[740])	,.Q4(Q[741])	,.Q5(Q[742])	,.Q6(Q[743])			,.R1(R[738])	,.R2(R[739])	,.R3(R[740])	,.R4(R[741])	,.R5(R[742])	,.R6(R[743])			,.clk(clk)	);
CNU_6 CNU117	(.Q1(Q[744])	,.Q2(Q[745])	,.Q3(Q[746])	,.Q4(Q[747])	,.Q5(Q[748])	,.Q6(Q[749])			,.R1(R[744])	,.R2(R[745])	,.R3(R[746])	,.R4(R[747])	,.R5(R[748])	,.R6(R[749])			,.clk(clk)	);
CNU_6 CNU118	(.Q1(Q[750])	,.Q2(Q[751])	,.Q3(Q[752])	,.Q4(Q[753])	,.Q5(Q[754])	,.Q6(Q[755])			,.R1(R[750])	,.R2(R[751])	,.R3(R[752])	,.R4(R[753])	,.R5(R[754])	,.R6(R[755])			,.clk(clk)	);
CNU_6 CNU119	(.Q1(Q[756])	,.Q2(Q[757])	,.Q3(Q[758])	,.Q4(Q[759])	,.Q5(Q[760])	,.Q6(Q[761])			,.R1(R[756])	,.R2(R[757])	,.R3(R[758])	,.R4(R[759])	,.R5(R[760])	,.R6(R[761])			,.clk(clk)	);
CNU_6 CNU120	(.Q1(Q[762])	,.Q2(Q[763])	,.Q3(Q[764])	,.Q4(Q[765])	,.Q5(Q[766])	,.Q6(Q[767])			,.R1(R[762])	,.R2(R[763])	,.R3(R[764])	,.R4(R[765])	,.R5(R[766])	,.R6(R[767])			,.clk(clk)	);

CNU_7 CNU121	(.Q1(Q[768])	,.Q2(Q[769])	,.Q3(Q[770])	,.Q4(Q[771])	,.Q5(Q[772])	,.Q6(Q[773])	,.Q7(Q[774])	,.R1(R[768])	,.R2(R[769])	,.R3(R[770])	,.R4(R[771])	,.R5(R[772])	,.R6(R[773])	,.R7(R[774])	,.clk(clk)	);
CNU_7 CNU122	(.Q1(Q[775])	,.Q2(Q[776])	,.Q3(Q[777])	,.Q4(Q[778])	,.Q5(Q[779])	,.Q6(Q[780])	,.Q7(Q[781])	,.R1(R[775])	,.R2(R[776])	,.R3(R[777])	,.R4(R[778])	,.R5(R[779])	,.R6(R[780])	,.R7(R[781])	,.clk(clk)	);
CNU_7 CNU123	(.Q1(Q[782])	,.Q2(Q[783])	,.Q3(Q[784])	,.Q4(Q[785])	,.Q5(Q[786])	,.Q6(Q[787])	,.Q7(Q[788])	,.R1(R[782])	,.R2(R[783])	,.R3(R[784])	,.R4(R[785])	,.R5(R[786])	,.R6(R[787])	,.R7(R[788])	,.clk(clk)	);
CNU_7 CNU124	(.Q1(Q[789])	,.Q2(Q[790])	,.Q3(Q[791])	,.Q4(Q[792])	,.Q5(Q[793])	,.Q6(Q[794])	,.Q7(Q[795])	,.R1(R[789])	,.R2(R[790])	,.R3(R[791])	,.R4(R[792])	,.R5(R[793])	,.R6(R[794])	,.R7(R[795])	,.clk(clk)	);
CNU_7 CNU125	(.Q1(Q[796])	,.Q2(Q[797])	,.Q3(Q[798])	,.Q4(Q[799])	,.Q5(Q[800])	,.Q6(Q[801])	,.Q7(Q[802])	,.R1(R[796])	,.R2(R[797])	,.R3(R[798])	,.R4(R[799])	,.R5(R[800])	,.R6(R[801])	,.R7(R[802])	,.clk(clk)	);
CNU_7 CNU126	(.Q1(Q[803])	,.Q2(Q[804])	,.Q3(Q[805])	,.Q4(Q[806])	,.Q5(Q[807])	,.Q6(Q[808])	,.Q7(Q[809])	,.R1(R[803])	,.R2(R[804])	,.R3(R[805])	,.R4(R[806])	,.R5(R[807])	,.R6(R[808])	,.R7(R[809])	,.clk(clk)	);
CNU_7 CNU127	(.Q1(Q[810])	,.Q2(Q[811])	,.Q3(Q[812])	,.Q4(Q[813])	,.Q5(Q[814])	,.Q6(Q[815])	,.Q7(Q[816])	,.R1(R[810])	,.R2(R[811])	,.R3(R[812])	,.R4(R[813])	,.R5(R[814])	,.R6(R[815])	,.R7(R[816])	,.clk(clk)	);
CNU_7 CNU128	(.Q1(Q[817])	,.Q2(Q[818])	,.Q3(Q[819])	,.Q4(Q[820])	,.Q5(Q[821])	,.Q6(Q[822])	,.Q7(Q[823])	,.R1(R[817])	,.R2(R[818])	,.R3(R[819])	,.R4(R[820])	,.R5(R[821])	,.R6(R[822])	,.R7(R[823])	,.clk(clk)	);
CNU_7 CNU129	(.Q1(Q[824])	,.Q2(Q[825])	,.Q3(Q[826])	,.Q4(Q[827])	,.Q5(Q[828])	,.Q6(Q[829])	,.Q7(Q[830])	,.R1(R[824])	,.R2(R[825])	,.R3(R[826])	,.R4(R[827])	,.R5(R[828])	,.R6(R[829])	,.R7(R[830])	,.clk(clk)	);
CNU_7 CNU130	(.Q1(Q[831])	,.Q2(Q[832])	,.Q3(Q[833])	,.Q4(Q[834])	,.Q5(Q[835])	,.Q6(Q[836])	,.Q7(Q[837])	,.R1(R[831])	,.R2(R[832])	,.R3(R[833])	,.R4(R[834])	,.R5(R[835])	,.R6(R[836])	,.R7(R[837])	,.clk(clk)	);
CNU_7 CNU131	(.Q1(Q[838])	,.Q2(Q[839])	,.Q3(Q[840])	,.Q4(Q[841])	,.Q5(Q[842])	,.Q6(Q[843])	,.Q7(Q[844])	,.R1(R[838])	,.R2(R[839])	,.R3(R[840])	,.R4(R[841])	,.R5(R[842])	,.R6(R[843])	,.R7(R[844])	,.clk(clk)	);
CNU_7 CNU132	(.Q1(Q[845])	,.Q2(Q[846])	,.Q3(Q[847])	,.Q4(Q[848])	,.Q5(Q[849])	,.Q6(Q[850])	,.Q7(Q[851])	,.R1(R[845])	,.R2(R[846])	,.R3(R[847])	,.R4(R[848])	,.R5(R[849])	,.R6(R[850])	,.R7(R[851])	,.clk(clk)	);
CNU_7 CNU133	(.Q1(Q[852])	,.Q2(Q[853])	,.Q3(Q[854])	,.Q4(Q[855])	,.Q5(Q[856])	,.Q6(Q[857])	,.Q7(Q[858])	,.R1(R[852])	,.R2(R[853])	,.R3(R[854])	,.R4(R[855])	,.R5(R[856])	,.R6(R[857])	,.R7(R[858])	,.clk(clk)	);
CNU_7 CNU134	(.Q1(Q[859])	,.Q2(Q[860])	,.Q3(Q[861])	,.Q4(Q[862])	,.Q5(Q[863])	,.Q6(Q[864])	,.Q7(Q[865])	,.R1(R[859])	,.R2(R[860])	,.R3(R[861])	,.R4(R[862])	,.R5(R[863])	,.R6(R[864])	,.R7(R[865])	,.clk(clk)	);
CNU_7 CNU135	(.Q1(Q[866])	,.Q2(Q[867])	,.Q3(Q[868])	,.Q4(Q[869])	,.Q5(Q[870])	,.Q6(Q[871])	,.Q7(Q[872])	,.R1(R[866])	,.R2(R[867])	,.R3(R[868])	,.R4(R[869])	,.R5(R[870])	,.R6(R[871])	,.R7(R[872])	,.clk(clk)	);
CNU_7 CNU136	(.Q1(Q[873])	,.Q2(Q[874])	,.Q3(Q[875])	,.Q4(Q[876])	,.Q5(Q[877])	,.Q6(Q[878])	,.Q7(Q[879])	,.R1(R[873])	,.R2(R[874])	,.R3(R[875])	,.R4(R[876])	,.R5(R[877])	,.R6(R[878])	,.R7(R[879])	,.clk(clk)	);
CNU_7 CNU137	(.Q1(Q[880])	,.Q2(Q[881])	,.Q3(Q[882])	,.Q4(Q[883])	,.Q5(Q[884])	,.Q6(Q[885])	,.Q7(Q[886])	,.R1(R[880])	,.R2(R[881])	,.R3(R[882])	,.R4(R[883])	,.R5(R[884])	,.R6(R[885])	,.R7(R[886])	,.clk(clk)	);
CNU_7 CNU138	(.Q1(Q[887])	,.Q2(Q[888])	,.Q3(Q[889])	,.Q4(Q[890])	,.Q5(Q[891])	,.Q6(Q[892])	,.Q7(Q[893])	,.R1(R[887])	,.R2(R[888])	,.R3(R[889])	,.R4(R[890])	,.R5(R[891])	,.R6(R[892])	,.R7(R[893])	,.clk(clk)	);
CNU_7 CNU139	(.Q1(Q[894])	,.Q2(Q[895])	,.Q3(Q[896])	,.Q4(Q[897])	,.Q5(Q[898])	,.Q6(Q[899])	,.Q7(Q[900])	,.R1(R[894])	,.R2(R[895])	,.R3(R[896])	,.R4(R[897])	,.R5(R[898])	,.R6(R[899])	,.R7(R[900])	,.clk(clk)	);
CNU_7 CNU140	(.Q1(Q[901])	,.Q2(Q[902])	,.Q3(Q[903])	,.Q4(Q[904])	,.Q5(Q[905])	,.Q6(Q[906])	,.Q7(Q[907])	,.R1(R[901])	,.R2(R[902])	,.R3(R[903])	,.R4(R[904])	,.R5(R[905])	,.R6(R[906])	,.R7(R[907])	,.clk(clk)	);
CNU_7 CNU141	(.Q1(Q[908])	,.Q2(Q[909])	,.Q3(Q[910])	,.Q4(Q[911])	,.Q5(Q[912])	,.Q6(Q[913])	,.Q7(Q[914])	,.R1(R[908])	,.R2(R[909])	,.R3(R[910])	,.R4(R[911])	,.R5(R[912])	,.R6(R[913])	,.R7(R[914])	,.clk(clk)	);
CNU_7 CNU142	(.Q1(Q[915])	,.Q2(Q[916])	,.Q3(Q[917])	,.Q4(Q[918])	,.Q5(Q[919])	,.Q6(Q[920])	,.Q7(Q[921])	,.R1(R[915])	,.R2(R[916])	,.R3(R[917])	,.R4(R[918])	,.R5(R[919])	,.R6(R[920])	,.R7(R[921])	,.clk(clk)	);
CNU_7 CNU143	(.Q1(Q[922])	,.Q2(Q[923])	,.Q3(Q[924])	,.Q4(Q[925])	,.Q5(Q[926])	,.Q6(Q[927])	,.Q7(Q[928])	,.R1(R[922])	,.R2(R[923])	,.R3(R[924])	,.R4(R[925])	,.R5(R[926])	,.R6(R[927])	,.R7(R[928])	,.clk(clk)	);
CNU_7 CNU144	(.Q1(Q[929])	,.Q2(Q[930])	,.Q3(Q[931])	,.Q4(Q[932])	,.Q5(Q[933])	,.Q6(Q[934])	,.Q7(Q[935])	,.R1(R[929])	,.R2(R[930])	,.R3(R[931])	,.R4(R[932])	,.R5(R[933])	,.R6(R[934])	,.R7(R[935])	,.clk(clk)	);

CNU_6 CNU145	(.Q1(Q[936])	,.Q2(Q[937])	,.Q3(Q[938])	,.Q4(Q[939])	,.Q5(Q[940])	,.Q6(Q[941])			,.R1(R[936])	,.R2(R[937])	,.R3(R[938])	,.R4(R[939])	,.R5(R[940])	,.R6(R[941])			,.clk(clk)	);
CNU_6 CNU146	(.Q1(Q[942])	,.Q2(Q[943])	,.Q3(Q[944])	,.Q4(Q[945])	,.Q5(Q[946])	,.Q6(Q[947])			,.R1(R[942])	,.R2(R[943])	,.R3(R[944])	,.R4(R[945])	,.R5(R[946])	,.R6(R[947])			,.clk(clk)	);
CNU_6 CNU147	(.Q1(Q[948])	,.Q2(Q[949])	,.Q3(Q[950])	,.Q4(Q[951])	,.Q5(Q[952])	,.Q6(Q[953])			,.R1(R[948])	,.R2(R[949])	,.R3(R[950])	,.R4(R[951])	,.R5(R[952])	,.R6(R[953])			,.clk(clk)	);
CNU_6 CNU148	(.Q1(Q[954])	,.Q2(Q[955])	,.Q3(Q[956])	,.Q4(Q[957])	,.Q5(Q[958])	,.Q6(Q[959])			,.R1(R[954])	,.R2(R[955])	,.R3(R[956])	,.R4(R[957])	,.R5(R[958])	,.R6(R[959])			,.clk(clk)	);
CNU_6 CNU149	(.Q1(Q[960])	,.Q2(Q[961])	,.Q3(Q[962])	,.Q4(Q[963])	,.Q5(Q[964])	,.Q6(Q[965])			,.R1(R[960])	,.R2(R[961])	,.R3(R[962])	,.R4(R[963])	,.R5(R[964])	,.R6(R[965])			,.clk(clk)	);
CNU_6 CNU150	(.Q1(Q[966])	,.Q2(Q[967])	,.Q3(Q[968])	,.Q4(Q[969])	,.Q5(Q[970])	,.Q6(Q[971])			,.R1(R[966])	,.R2(R[967])	,.R3(R[968])	,.R4(R[969])	,.R5(R[970])	,.R6(R[971])			,.clk(clk)	);
CNU_6 CNU151	(.Q1(Q[972])	,.Q2(Q[973])	,.Q3(Q[974])	,.Q4(Q[975])	,.Q5(Q[976])	,.Q6(Q[977])			,.R1(R[972])	,.R2(R[973])	,.R3(R[974])	,.R4(R[975])	,.R5(R[976])	,.R6(R[977])			,.clk(clk)	);
CNU_6 CNU152	(.Q1(Q[978])	,.Q2(Q[979])	,.Q3(Q[980])	,.Q4(Q[981])	,.Q5(Q[982])	,.Q6(Q[983])			,.R1(R[978])	,.R2(R[979])	,.R3(R[980])	,.R4(R[981])	,.R5(R[982])	,.R6(R[983])			,.clk(clk)	);
CNU_6 CNU153	(.Q1(Q[984])	,.Q2(Q[985])	,.Q3(Q[986])	,.Q4(Q[987])	,.Q5(Q[988])	,.Q6(Q[989])			,.R1(R[984])	,.R2(R[985])	,.R3(R[986])	,.R4(R[987])	,.R5(R[988])	,.R6(R[989])			,.clk(clk)	);
CNU_6 CNU154	(.Q1(Q[990])	,.Q2(Q[991])	,.Q3(Q[992])	,.Q4(Q[993])	,.Q5(Q[994])	,.Q6(Q[995])			,.R1(R[990])	,.R2(R[991])	,.R3(R[992])	,.R4(R[993])	,.R5(R[994])	,.R6(R[995])			,.clk(clk)	);
CNU_6 CNU155	(.Q1(Q[996])	,.Q2(Q[997])	,.Q3(Q[998])	,.Q4(Q[999])	,.Q5(Q[1000])	,.Q6(Q[1001])			,.R1(R[996])	,.R2(R[997])	,.R3(R[998])	,.R4(R[999])	,.R5(R[1000])	,.R6(R[1001])			,.clk(clk)	);
CNU_6 CNU156	(.Q1(Q[1002])	,.Q2(Q[1003])	,.Q3(Q[1004])	,.Q4(Q[1005])	,.Q5(Q[1006])	,.Q6(Q[1007])			,.R1(R[1002])	,.R2(R[1003])	,.R3(R[1004])	,.R4(R[1005])	,.R5(R[1006])	,.R6(R[1007])			,.clk(clk)	);
CNU_6 CNU157	(.Q1(Q[1008])	,.Q2(Q[1009])	,.Q3(Q[1010])	,.Q4(Q[1011])	,.Q5(Q[1012])	,.Q6(Q[1013])			,.R1(R[1008])	,.R2(R[1009])	,.R3(R[1010])	,.R4(R[1011])	,.R5(R[1012])	,.R6(R[1013])			,.clk(clk)	);
CNU_6 CNU158	(.Q1(Q[1014])	,.Q2(Q[1015])	,.Q3(Q[1016])	,.Q4(Q[1017])	,.Q5(Q[1018])	,.Q6(Q[1019])			,.R1(R[1014])	,.R2(R[1015])	,.R3(R[1016])	,.R4(R[1017])	,.R5(R[1018])	,.R6(R[1019])			,.clk(clk)	);
CNU_6 CNU159	(.Q1(Q[1020])	,.Q2(Q[1021])	,.Q3(Q[1022])	,.Q4(Q[1023])	,.Q5(Q[1024])	,.Q6(Q[1025])			,.R1(R[1020])	,.R2(R[1021])	,.R3(R[1022])	,.R4(R[1023])	,.R5(R[1024])	,.R6(R[1025])			,.clk(clk)	);
CNU_6 CNU160	(.Q1(Q[1026])	,.Q2(Q[1027])	,.Q3(Q[1028])	,.Q4(Q[1029])	,.Q5(Q[1030])	,.Q6(Q[1031])			,.R1(R[1026])	,.R2(R[1027])	,.R3(R[1028])	,.R4(R[1029])	,.R5(R[1030])	,.R6(R[1031])			,.clk(clk)	);
CNU_6 CNU161	(.Q1(Q[1032])	,.Q2(Q[1033])	,.Q3(Q[1034])	,.Q4(Q[1035])	,.Q5(Q[1036])	,.Q6(Q[1037])			,.R1(R[1032])	,.R2(R[1033])	,.R3(R[1034])	,.R4(R[1035])	,.R5(R[1036])	,.R6(R[1037])			,.clk(clk)	);
CNU_6 CNU162	(.Q1(Q[1038])	,.Q2(Q[1039])	,.Q3(Q[1040])	,.Q4(Q[1041])	,.Q5(Q[1042])	,.Q6(Q[1043])			,.R1(R[1038])	,.R2(R[1039])	,.R3(R[1040])	,.R4(R[1041])	,.R5(R[1042])	,.R6(R[1043])			,.clk(clk)	);
CNU_6 CNU163	(.Q1(Q[1044])	,.Q2(Q[1045])	,.Q3(Q[1046])	,.Q4(Q[1047])	,.Q5(Q[1048])	,.Q6(Q[1049])			,.R1(R[1044])	,.R2(R[1045])	,.R3(R[1046])	,.R4(R[1047])	,.R5(R[1048])	,.R6(R[1049])			,.clk(clk)	);
CNU_6 CNU164	(.Q1(Q[1050])	,.Q2(Q[1051])	,.Q3(Q[1052])	,.Q4(Q[1053])	,.Q5(Q[1054])	,.Q6(Q[1055])			,.R1(R[1050])	,.R2(R[1051])	,.R3(R[1052])	,.R4(R[1053])	,.R5(R[1054])	,.R6(R[1055])			,.clk(clk)	);
CNU_6 CNU165	(.Q1(Q[1056])	,.Q2(Q[1057])	,.Q3(Q[1058])	,.Q4(Q[1059])	,.Q5(Q[1060])	,.Q6(Q[1061])			,.R1(R[1056])	,.R2(R[1057])	,.R3(R[1058])	,.R4(R[1059])	,.R5(R[1060])	,.R6(R[1061])			,.clk(clk)	);
CNU_6 CNU166	(.Q1(Q[1062])	,.Q2(Q[1063])	,.Q3(Q[1064])	,.Q4(Q[1065])	,.Q5(Q[1066])	,.Q6(Q[1067])			,.R1(R[1062])	,.R2(R[1063])	,.R3(R[1064])	,.R4(R[1065])	,.R5(R[1066])	,.R6(R[1067])			,.clk(clk)	);
CNU_6 CNU167	(.Q1(Q[1068])	,.Q2(Q[1069])	,.Q3(Q[1070])	,.Q4(Q[1071])	,.Q5(Q[1072])	,.Q6(Q[1073])			,.R1(R[1068])	,.R2(R[1069])	,.R3(R[1070])	,.R4(R[1071])	,.R5(R[1072])	,.R6(R[1073])			,.clk(clk)	);
CNU_6 CNU168	(.Q1(Q[1074])	,.Q2(Q[1075])	,.Q3(Q[1076])	,.Q4(Q[1077])	,.Q5(Q[1078])	,.Q6(Q[1079])			,.R1(R[1074])	,.R2(R[1075])	,.R3(R[1076])	,.R4(R[1077])	,.R5(R[1078])	,.R6(R[1079])			,.clk(clk)	);
CNU_6 CNU169	(.Q1(Q[1080])	,.Q2(Q[1081])	,.Q3(Q[1082])	,.Q4(Q[1083])	,.Q5(Q[1084])	,.Q6(Q[1085])			,.R1(R[1080])	,.R2(R[1081])	,.R3(R[1082])	,.R4(R[1083])	,.R5(R[1084])	,.R6(R[1085])			,.clk(clk)	);
CNU_6 CNU170	(.Q1(Q[1086])	,.Q2(Q[1087])	,.Q3(Q[1088])	,.Q4(Q[1089])	,.Q5(Q[1090])	,.Q6(Q[1091])			,.R1(R[1086])	,.R2(R[1087])	,.R3(R[1088])	,.R4(R[1089])	,.R5(R[1090])	,.R6(R[1091])			,.clk(clk)	);
CNU_6 CNU171	(.Q1(Q[1092])	,.Q2(Q[1093])	,.Q3(Q[1094])	,.Q4(Q[1095])	,.Q5(Q[1096])	,.Q6(Q[1097])			,.R1(R[1092])	,.R2(R[1093])	,.R3(R[1094])	,.R4(R[1095])	,.R5(R[1096])	,.R6(R[1097])			,.clk(clk)	);
CNU_6 CNU172	(.Q1(Q[1098])	,.Q2(Q[1099])	,.Q3(Q[1100])	,.Q4(Q[1101])	,.Q5(Q[1102])	,.Q6(Q[1103])			,.R1(R[1098])	,.R2(R[1099])	,.R3(R[1100])	,.R4(R[1101])	,.R5(R[1102])	,.R6(R[1103])			,.clk(clk)	);
CNU_6 CNU173	(.Q1(Q[1104])	,.Q2(Q[1105])	,.Q3(Q[1106])	,.Q4(Q[1107])	,.Q5(Q[1108])	,.Q6(Q[1109])			,.R1(R[1104])	,.R2(R[1105])	,.R3(R[1106])	,.R4(R[1107])	,.R5(R[1108])	,.R6(R[1109])			,.clk(clk)	);
CNU_6 CNU174	(.Q1(Q[1110])	,.Q2(Q[1111])	,.Q3(Q[1112])	,.Q4(Q[1113])	,.Q5(Q[1114])	,.Q6(Q[1115])			,.R1(R[1110])	,.R2(R[1111])	,.R3(R[1112])	,.R4(R[1113])	,.R5(R[1114])	,.R6(R[1115])			,.clk(clk)	);
CNU_6 CNU175	(.Q1(Q[1116])	,.Q2(Q[1117])	,.Q3(Q[1118])	,.Q4(Q[1119])	,.Q5(Q[1120])	,.Q6(Q[1121])			,.R1(R[1116])	,.R2(R[1117])	,.R3(R[1118])	,.R4(R[1119])	,.R5(R[1120])	,.R6(R[1121])			,.clk(clk)	);
CNU_6 CNU176	(.Q1(Q[1122])	,.Q2(Q[1123])	,.Q3(Q[1124])	,.Q4(Q[1125])	,.Q5(Q[1126])	,.Q6(Q[1127])			,.R1(R[1122])	,.R2(R[1123])	,.R3(R[1124])	,.R4(R[1125])	,.R5(R[1126])	,.R6(R[1127])			,.clk(clk)	);
CNU_6 CNU177	(.Q1(Q[1128])	,.Q2(Q[1129])	,.Q3(Q[1130])	,.Q4(Q[1131])	,.Q5(Q[1132])	,.Q6(Q[1133])			,.R1(R[1128])	,.R2(R[1129])	,.R3(R[1130])	,.R4(R[1131])	,.R5(R[1132])	,.R6(R[1133])			,.clk(clk)	);
CNU_6 CNU178	(.Q1(Q[1134])	,.Q2(Q[1135])	,.Q3(Q[1136])	,.Q4(Q[1137])	,.Q5(Q[1138])	,.Q6(Q[1139])			,.R1(R[1134])	,.R2(R[1135])	,.R3(R[1136])	,.R4(R[1137])	,.R5(R[1138])	,.R6(R[1139])			,.clk(clk)	);
CNU_6 CNU179	(.Q1(Q[1140])	,.Q2(Q[1141])	,.Q3(Q[1142])	,.Q4(Q[1143])	,.Q5(Q[1144])	,.Q6(Q[1145])			,.R1(R[1140])	,.R2(R[1141])	,.R3(R[1142])	,.R4(R[1143])	,.R5(R[1144])	,.R6(R[1145])			,.clk(clk)	);
CNU_6 CNU180	(.Q1(Q[1146])	,.Q2(Q[1147])	,.Q3(Q[1148])	,.Q4(Q[1149])	,.Q5(Q[1150])	,.Q6(Q[1151])			,.R1(R[1146])	,.R2(R[1147])	,.R3(R[1148])	,.R4(R[1149])	,.R5(R[1150])	,.R6(R[1151])			,.clk(clk)	);
CNU_6 CNU181	(.Q1(Q[1152])	,.Q2(Q[1153])	,.Q3(Q[1154])	,.Q4(Q[1155])	,.Q5(Q[1156])	,.Q6(Q[1157])			,.R1(R[1152])	,.R2(R[1153])	,.R3(R[1154])	,.R4(R[1155])	,.R5(R[1156])	,.R6(R[1157])			,.clk(clk)	);
CNU_6 CNU182	(.Q1(Q[1158])	,.Q2(Q[1159])	,.Q3(Q[1160])	,.Q4(Q[1161])	,.Q5(Q[1162])	,.Q6(Q[1163])			,.R1(R[1158])	,.R2(R[1159])	,.R3(R[1160])	,.R4(R[1161])	,.R5(R[1162])	,.R6(R[1163])			,.clk(clk)	);
CNU_6 CNU183	(.Q1(Q[1164])	,.Q2(Q[1165])	,.Q3(Q[1166])	,.Q4(Q[1167])	,.Q5(Q[1168])	,.Q6(Q[1169])			,.R1(R[1164])	,.R2(R[1165])	,.R3(R[1166])	,.R4(R[1167])	,.R5(R[1168])	,.R6(R[1169])			,.clk(clk)	);
CNU_6 CNU184	(.Q1(Q[1170])	,.Q2(Q[1171])	,.Q3(Q[1172])	,.Q4(Q[1173])	,.Q5(Q[1174])	,.Q6(Q[1175])			,.R1(R[1170])	,.R2(R[1171])	,.R3(R[1172])	,.R4(R[1173])	,.R5(R[1174])	,.R6(R[1175])			,.clk(clk)	);
CNU_6 CNU185	(.Q1(Q[1176])	,.Q2(Q[1177])	,.Q3(Q[1178])	,.Q4(Q[1179])	,.Q5(Q[1180])	,.Q6(Q[1181])			,.R1(R[1176])	,.R2(R[1177])	,.R3(R[1178])	,.R4(R[1179])	,.R5(R[1180])	,.R6(R[1181])			,.clk(clk)	);
CNU_6 CNU186	(.Q1(Q[1182])	,.Q2(Q[1183])	,.Q3(Q[1184])	,.Q4(Q[1185])	,.Q5(Q[1186])	,.Q6(Q[1187])			,.R1(R[1182])	,.R2(R[1183])	,.R3(R[1184])	,.R4(R[1185])	,.R5(R[1186])	,.R6(R[1187])			,.clk(clk)	);
CNU_6 CNU187	(.Q1(Q[1188])	,.Q2(Q[1189])	,.Q3(Q[1190])	,.Q4(Q[1191])	,.Q5(Q[1192])	,.Q6(Q[1193])			,.R1(R[1188])	,.R2(R[1189])	,.R3(R[1190])	,.R4(R[1191])	,.R5(R[1192])	,.R6(R[1193])			,.clk(clk)	);
CNU_6 CNU188	(.Q1(Q[1194])	,.Q2(Q[1195])	,.Q3(Q[1196])	,.Q4(Q[1197])	,.Q5(Q[1198])	,.Q6(Q[1199])			,.R1(R[1194])	,.R2(R[1195])	,.R3(R[1196])	,.R4(R[1197])	,.R5(R[1198])	,.R6(R[1199])			,.clk(clk)	);
CNU_6 CNU189	(.Q1(Q[1200])	,.Q2(Q[1201])	,.Q3(Q[1202])	,.Q4(Q[1203])	,.Q5(Q[1204])	,.Q6(Q[1205])			,.R1(R[1200])	,.R2(R[1201])	,.R3(R[1202])	,.R4(R[1203])	,.R5(R[1204])	,.R6(R[1205])			,.clk(clk)	);
CNU_6 CNU190	(.Q1(Q[1206])	,.Q2(Q[1207])	,.Q3(Q[1208])	,.Q4(Q[1209])	,.Q5(Q[1210])	,.Q6(Q[1211])			,.R1(R[1206])	,.R2(R[1207])	,.R3(R[1208])	,.R4(R[1209])	,.R5(R[1210])	,.R6(R[1211])			,.clk(clk)	);
CNU_6 CNU191	(.Q1(Q[1212])	,.Q2(Q[1213])	,.Q3(Q[1214])	,.Q4(Q[1215])	,.Q5(Q[1216])	,.Q6(Q[1217])			,.R1(R[1212])	,.R2(R[1213])	,.R3(R[1214])	,.R4(R[1215])	,.R5(R[1216])	,.R6(R[1217])			,.clk(clk)	);
CNU_6 CNU192	(.Q1(Q[1218])	,.Q2(Q[1219])	,.Q3(Q[1220])	,.Q4(Q[1221])	,.Q5(Q[1222])	,.Q6(Q[1223])			,.R1(R[1218])	,.R2(R[1219])	,.R3(R[1220])	,.R4(R[1221])	,.R5(R[1222])	,.R6(R[1223])			,.clk(clk)	);

CNU_7 CNU193	(.Q1(Q[1224])	,.Q2(Q[1225])	,.Q3(Q[1226])	,.Q4(Q[1227])	,.Q5(Q[1228])	,.Q6(Q[1229])	,.Q7(Q[1230])	,.R1(R[1224])	,.R2(R[1225])	,.R3(R[1226])	,.R4(R[1227])	,.R5(R[1228])	,.R6(R[1229])	,.R7(R[1230])	,.clk(clk)	);
CNU_7 CNU194	(.Q1(Q[1231])	,.Q2(Q[1232])	,.Q3(Q[1233])	,.Q4(Q[1234])	,.Q5(Q[1235])	,.Q6(Q[1236])	,.Q7(Q[1237])	,.R1(R[1231])	,.R2(R[1232])	,.R3(R[1233])	,.R4(R[1234])	,.R5(R[1235])	,.R6(R[1236])	,.R7(R[1237])	,.clk(clk)	);
CNU_7 CNU195	(.Q1(Q[1238])	,.Q2(Q[1239])	,.Q3(Q[1240])	,.Q4(Q[1241])	,.Q5(Q[1242])	,.Q6(Q[1243])	,.Q7(Q[1244])	,.R1(R[1238])	,.R2(R[1239])	,.R3(R[1240])	,.R4(R[1241])	,.R5(R[1242])	,.R6(R[1243])	,.R7(R[1244])	,.clk(clk)	);
CNU_7 CNU196	(.Q1(Q[1245])	,.Q2(Q[1246])	,.Q3(Q[1247])	,.Q4(Q[1248])	,.Q5(Q[1249])	,.Q6(Q[1250])	,.Q7(Q[1251])	,.R1(R[1245])	,.R2(R[1246])	,.R3(R[1247])	,.R4(R[1248])	,.R5(R[1249])	,.R6(R[1250])	,.R7(R[1251])	,.clk(clk)	);
CNU_7 CNU197	(.Q1(Q[1252])	,.Q2(Q[1253])	,.Q3(Q[1254])	,.Q4(Q[1255])	,.Q5(Q[1256])	,.Q6(Q[1257])	,.Q7(Q[1258])	,.R1(R[1252])	,.R2(R[1253])	,.R3(R[1254])	,.R4(R[1255])	,.R5(R[1256])	,.R6(R[1257])	,.R7(R[1258])	,.clk(clk)	);
CNU_7 CNU198	(.Q1(Q[1259])	,.Q2(Q[1260])	,.Q3(Q[1261])	,.Q4(Q[1262])	,.Q5(Q[1263])	,.Q6(Q[1264])	,.Q7(Q[1265])	,.R1(R[1259])	,.R2(R[1260])	,.R3(R[1261])	,.R4(R[1262])	,.R5(R[1263])	,.R6(R[1264])	,.R7(R[1265])	,.clk(clk)	);
CNU_7 CNU199	(.Q1(Q[1266])	,.Q2(Q[1267])	,.Q3(Q[1268])	,.Q4(Q[1269])	,.Q5(Q[1270])	,.Q6(Q[1271])	,.Q7(Q[1272])	,.R1(R[1266])	,.R2(R[1267])	,.R3(R[1268])	,.R4(R[1269])	,.R5(R[1270])	,.R6(R[1271])	,.R7(R[1272])	,.clk(clk)	);
CNU_7 CNU200	(.Q1(Q[1273])	,.Q2(Q[1274])	,.Q3(Q[1275])	,.Q4(Q[1276])	,.Q5(Q[1277])	,.Q6(Q[1278])	,.Q7(Q[1279])	,.R1(R[1273])	,.R2(R[1274])	,.R3(R[1275])	,.R4(R[1276])	,.R5(R[1277])	,.R6(R[1278])	,.R7(R[1279])	,.clk(clk)	);
CNU_7 CNU201	(.Q1(Q[1280])	,.Q2(Q[1281])	,.Q3(Q[1282])	,.Q4(Q[1283])	,.Q5(Q[1284])	,.Q6(Q[1285])	,.Q7(Q[1286])	,.R1(R[1280])	,.R2(R[1281])	,.R3(R[1282])	,.R4(R[1283])	,.R5(R[1284])	,.R6(R[1285])	,.R7(R[1286])	,.clk(clk)	);
CNU_7 CNU202	(.Q1(Q[1287])	,.Q2(Q[1288])	,.Q3(Q[1289])	,.Q4(Q[1290])	,.Q5(Q[1291])	,.Q6(Q[1292])	,.Q7(Q[1293])	,.R1(R[1287])	,.R2(R[1288])	,.R3(R[1289])	,.R4(R[1290])	,.R5(R[1291])	,.R6(R[1292])	,.R7(R[1293])	,.clk(clk)	);
CNU_7 CNU203	(.Q1(Q[1294])	,.Q2(Q[1295])	,.Q3(Q[1296])	,.Q4(Q[1297])	,.Q5(Q[1298])	,.Q6(Q[1299])	,.Q7(Q[1300])	,.R1(R[1294])	,.R2(R[1295])	,.R3(R[1296])	,.R4(R[1297])	,.R5(R[1298])	,.R6(R[1299])	,.R7(R[1300])	,.clk(clk)	);
CNU_7 CNU204	(.Q1(Q[1301])	,.Q2(Q[1302])	,.Q3(Q[1303])	,.Q4(Q[1304])	,.Q5(Q[1305])	,.Q6(Q[1306])	,.Q7(Q[1307])	,.R1(R[1301])	,.R2(R[1302])	,.R3(R[1303])	,.R4(R[1304])	,.R5(R[1305])	,.R6(R[1306])	,.R7(R[1307])	,.clk(clk)	);
CNU_7 CNU205	(.Q1(Q[1308])	,.Q2(Q[1309])	,.Q3(Q[1310])	,.Q4(Q[1311])	,.Q5(Q[1312])	,.Q6(Q[1313])	,.Q7(Q[1314])	,.R1(R[1308])	,.R2(R[1309])	,.R3(R[1310])	,.R4(R[1311])	,.R5(R[1312])	,.R6(R[1313])	,.R7(R[1314])	,.clk(clk)	);
CNU_7 CNU206	(.Q1(Q[1315])	,.Q2(Q[1316])	,.Q3(Q[1317])	,.Q4(Q[1318])	,.Q5(Q[1319])	,.Q6(Q[1320])	,.Q7(Q[1321])	,.R1(R[1315])	,.R2(R[1316])	,.R3(R[1317])	,.R4(R[1318])	,.R5(R[1319])	,.R6(R[1320])	,.R7(R[1321])	,.clk(clk)	);
CNU_7 CNU207	(.Q1(Q[1322])	,.Q2(Q[1323])	,.Q3(Q[1324])	,.Q4(Q[1325])	,.Q5(Q[1326])	,.Q6(Q[1327])	,.Q7(Q[1328])	,.R1(R[1322])	,.R2(R[1323])	,.R3(R[1324])	,.R4(R[1325])	,.R5(R[1326])	,.R6(R[1327])	,.R7(R[1328])	,.clk(clk)	);
CNU_7 CNU208	(.Q1(Q[1329])	,.Q2(Q[1330])	,.Q3(Q[1331])	,.Q4(Q[1332])	,.Q5(Q[1333])	,.Q6(Q[1334])	,.Q7(Q[1335])	,.R1(R[1329])	,.R2(R[1330])	,.R3(R[1331])	,.R4(R[1332])	,.R5(R[1333])	,.R6(R[1334])	,.R7(R[1335])	,.clk(clk)	);
CNU_7 CNU209	(.Q1(Q[1336])	,.Q2(Q[1337])	,.Q3(Q[1338])	,.Q4(Q[1339])	,.Q5(Q[1340])	,.Q6(Q[1341])	,.Q7(Q[1342])	,.R1(R[1336])	,.R2(R[1337])	,.R3(R[1338])	,.R4(R[1339])	,.R5(R[1340])	,.R6(R[1341])	,.R7(R[1342])	,.clk(clk)	);
CNU_7 CNU210	(.Q1(Q[1343])	,.Q2(Q[1344])	,.Q3(Q[1345])	,.Q4(Q[1346])	,.Q5(Q[1347])	,.Q6(Q[1348])	,.Q7(Q[1349])	,.R1(R[1343])	,.R2(R[1344])	,.R3(R[1345])	,.R4(R[1346])	,.R5(R[1347])	,.R6(R[1348])	,.R7(R[1349])	,.clk(clk)	);
CNU_7 CNU211	(.Q1(Q[1350])	,.Q2(Q[1351])	,.Q3(Q[1352])	,.Q4(Q[1353])	,.Q5(Q[1354])	,.Q6(Q[1355])	,.Q7(Q[1356])	,.R1(R[1350])	,.R2(R[1351])	,.R3(R[1352])	,.R4(R[1353])	,.R5(R[1354])	,.R6(R[1355])	,.R7(R[1356])	,.clk(clk)	);
CNU_7 CNU212	(.Q1(Q[1357])	,.Q2(Q[1358])	,.Q3(Q[1359])	,.Q4(Q[1360])	,.Q5(Q[1361])	,.Q6(Q[1362])	,.Q7(Q[1363])	,.R1(R[1357])	,.R2(R[1358])	,.R3(R[1359])	,.R4(R[1360])	,.R5(R[1361])	,.R6(R[1362])	,.R7(R[1363])	,.clk(clk)	);
CNU_7 CNU213	(.Q1(Q[1364])	,.Q2(Q[1365])	,.Q3(Q[1366])	,.Q4(Q[1367])	,.Q5(Q[1368])	,.Q6(Q[1369])	,.Q7(Q[1370])	,.R1(R[1364])	,.R2(R[1365])	,.R3(R[1366])	,.R4(R[1367])	,.R5(R[1368])	,.R6(R[1369])	,.R7(R[1370])	,.clk(clk)	);
CNU_7 CNU214	(.Q1(Q[1371])	,.Q2(Q[1372])	,.Q3(Q[1373])	,.Q4(Q[1374])	,.Q5(Q[1375])	,.Q6(Q[1376])	,.Q7(Q[1377])	,.R1(R[1371])	,.R2(R[1372])	,.R3(R[1373])	,.R4(R[1374])	,.R5(R[1375])	,.R6(R[1376])	,.R7(R[1377])	,.clk(clk)	);
CNU_7 CNU215	(.Q1(Q[1378])	,.Q2(Q[1379])	,.Q3(Q[1380])	,.Q4(Q[1381])	,.Q5(Q[1382])	,.Q6(Q[1383])	,.Q7(Q[1384])	,.R1(R[1378])	,.R2(R[1379])	,.R3(R[1380])	,.R4(R[1381])	,.R5(R[1382])	,.R6(R[1383])	,.R7(R[1384])	,.clk(clk)	);
CNU_7 CNU216	(.Q1(Q[1385])	,.Q2(Q[1386])	,.Q3(Q[1387])	,.Q4(Q[1388])	,.Q5(Q[1389])	,.Q6(Q[1390])	,.Q7(Q[1391])	,.R1(R[1385])	,.R2(R[1386])	,.R3(R[1387])	,.R4(R[1388])	,.R5(R[1389])	,.R6(R[1390])	,.R7(R[1391])	,.clk(clk)	);

CNU_6 CNU217	(.Q1(Q[1392])	,.Q2(Q[1393])	,.Q3(Q[1394])	,.Q4(Q[1395])	,.Q5(Q[1396])	,.Q6(Q[1397])			,.R1(R[1392])	,.R2(R[1393])	,.R3(R[1394])	,.R4(R[1395])	,.R5(R[1396])	,.R6(R[1397])			,.clk(clk)	);
CNU_6 CNU218	(.Q1(Q[1398])	,.Q2(Q[1399])	,.Q3(Q[1400])	,.Q4(Q[1401])	,.Q5(Q[1402])	,.Q6(Q[1403])			,.R1(R[1398])	,.R2(R[1399])	,.R3(R[1400])	,.R4(R[1401])	,.R5(R[1402])	,.R6(R[1403])			,.clk(clk)	);
CNU_6 CNU219	(.Q1(Q[1404])	,.Q2(Q[1405])	,.Q3(Q[1406])	,.Q4(Q[1407])	,.Q5(Q[1408])	,.Q6(Q[1409])			,.R1(R[1404])	,.R2(R[1405])	,.R3(R[1406])	,.R4(R[1407])	,.R5(R[1408])	,.R6(R[1409])			,.clk(clk)	);
CNU_6 CNU220	(.Q1(Q[1410])	,.Q2(Q[1411])	,.Q3(Q[1412])	,.Q4(Q[1413])	,.Q5(Q[1414])	,.Q6(Q[1415])			,.R1(R[1410])	,.R2(R[1411])	,.R3(R[1412])	,.R4(R[1413])	,.R5(R[1414])	,.R6(R[1415])			,.clk(clk)	);
CNU_6 CNU221	(.Q1(Q[1416])	,.Q2(Q[1417])	,.Q3(Q[1418])	,.Q4(Q[1419])	,.Q5(Q[1420])	,.Q6(Q[1421])			,.R1(R[1416])	,.R2(R[1417])	,.R3(R[1418])	,.R4(R[1419])	,.R5(R[1420])	,.R6(R[1421])			,.clk(clk)	);
CNU_6 CNU222	(.Q1(Q[1422])	,.Q2(Q[1423])	,.Q3(Q[1424])	,.Q4(Q[1425])	,.Q5(Q[1426])	,.Q6(Q[1427])			,.R1(R[1422])	,.R2(R[1423])	,.R3(R[1424])	,.R4(R[1425])	,.R5(R[1426])	,.R6(R[1427])			,.clk(clk)	);
CNU_6 CNU223	(.Q1(Q[1428])	,.Q2(Q[1429])	,.Q3(Q[1430])	,.Q4(Q[1431])	,.Q5(Q[1432])	,.Q6(Q[1433])			,.R1(R[1428])	,.R2(R[1429])	,.R3(R[1430])	,.R4(R[1431])	,.R5(R[1432])	,.R6(R[1433])			,.clk(clk)	);
CNU_6 CNU224	(.Q1(Q[1434])	,.Q2(Q[1435])	,.Q3(Q[1436])	,.Q4(Q[1437])	,.Q5(Q[1438])	,.Q6(Q[1439])			,.R1(R[1434])	,.R2(R[1435])	,.R3(R[1436])	,.R4(R[1437])	,.R5(R[1438])	,.R6(R[1439])			,.clk(clk)	);
CNU_6 CNU225	(.Q1(Q[1440])	,.Q2(Q[1441])	,.Q3(Q[1442])	,.Q4(Q[1443])	,.Q5(Q[1444])	,.Q6(Q[1445])			,.R1(R[1440])	,.R2(R[1441])	,.R3(R[1442])	,.R4(R[1443])	,.R5(R[1444])	,.R6(R[1445])			,.clk(clk)	);
CNU_6 CNU226	(.Q1(Q[1446])	,.Q2(Q[1447])	,.Q3(Q[1448])	,.Q4(Q[1449])	,.Q5(Q[1450])	,.Q6(Q[1451])			,.R1(R[1446])	,.R2(R[1447])	,.R3(R[1448])	,.R4(R[1449])	,.R5(R[1450])	,.R6(R[1451])			,.clk(clk)	);
CNU_6 CNU227	(.Q1(Q[1452])	,.Q2(Q[1453])	,.Q3(Q[1454])	,.Q4(Q[1455])	,.Q5(Q[1456])	,.Q6(Q[1457])			,.R1(R[1452])	,.R2(R[1453])	,.R3(R[1454])	,.R4(R[1455])	,.R5(R[1456])	,.R6(R[1457])			,.clk(clk)	);
CNU_6 CNU228	(.Q1(Q[1458])	,.Q2(Q[1459])	,.Q3(Q[1460])	,.Q4(Q[1461])	,.Q5(Q[1462])	,.Q6(Q[1463])			,.R1(R[1458])	,.R2(R[1459])	,.R3(R[1460])	,.R4(R[1461])	,.R5(R[1462])	,.R6(R[1463])			,.clk(clk)	);
CNU_6 CNU229	(.Q1(Q[1464])	,.Q2(Q[1465])	,.Q3(Q[1466])	,.Q4(Q[1467])	,.Q5(Q[1468])	,.Q6(Q[1469])			,.R1(R[1464])	,.R2(R[1465])	,.R3(R[1466])	,.R4(R[1467])	,.R5(R[1468])	,.R6(R[1469])			,.clk(clk)	);
CNU_6 CNU230	(.Q1(Q[1470])	,.Q2(Q[1471])	,.Q3(Q[1472])	,.Q4(Q[1473])	,.Q5(Q[1474])	,.Q6(Q[1475])			,.R1(R[1470])	,.R2(R[1471])	,.R3(R[1472])	,.R4(R[1473])	,.R5(R[1474])	,.R6(R[1475])			,.clk(clk)	);
CNU_6 CNU231	(.Q1(Q[1476])	,.Q2(Q[1477])	,.Q3(Q[1478])	,.Q4(Q[1479])	,.Q5(Q[1480])	,.Q6(Q[1481])			,.R1(R[1476])	,.R2(R[1477])	,.R3(R[1478])	,.R4(R[1479])	,.R5(R[1480])	,.R6(R[1481])			,.clk(clk)	);
CNU_6 CNU232	(.Q1(Q[1482])	,.Q2(Q[1483])	,.Q3(Q[1484])	,.Q4(Q[1485])	,.Q5(Q[1486])	,.Q6(Q[1487])			,.R1(R[1482])	,.R2(R[1483])	,.R3(R[1484])	,.R4(R[1485])	,.R5(R[1486])	,.R6(R[1487])			,.clk(clk)	);
CNU_6 CNU233	(.Q1(Q[1488])	,.Q2(Q[1489])	,.Q3(Q[1490])	,.Q4(Q[1491])	,.Q5(Q[1492])	,.Q6(Q[1493])			,.R1(R[1488])	,.R2(R[1489])	,.R3(R[1490])	,.R4(R[1491])	,.R5(R[1492])	,.R6(R[1493])			,.clk(clk)	);
CNU_6 CNU234	(.Q1(Q[1494])	,.Q2(Q[1495])	,.Q3(Q[1496])	,.Q4(Q[1497])	,.Q5(Q[1498])	,.Q6(Q[1499])			,.R1(R[1494])	,.R2(R[1495])	,.R3(R[1496])	,.R4(R[1497])	,.R5(R[1498])	,.R6(R[1499])			,.clk(clk)	);
CNU_6 CNU235	(.Q1(Q[1500])	,.Q2(Q[1501])	,.Q3(Q[1502])	,.Q4(Q[1503])	,.Q5(Q[1504])	,.Q6(Q[1505])			,.R1(R[1500])	,.R2(R[1501])	,.R3(R[1502])	,.R4(R[1503])	,.R5(R[1504])	,.R6(R[1505])			,.clk(clk)	);
CNU_6 CNU236	(.Q1(Q[1506])	,.Q2(Q[1507])	,.Q3(Q[1508])	,.Q4(Q[1509])	,.Q5(Q[1510])	,.Q6(Q[1511])			,.R1(R[1506])	,.R2(R[1507])	,.R3(R[1508])	,.R4(R[1509])	,.R5(R[1510])	,.R6(R[1511])			,.clk(clk)	);
CNU_6 CNU237	(.Q1(Q[1512])	,.Q2(Q[1513])	,.Q3(Q[1514])	,.Q4(Q[1515])	,.Q5(Q[1516])	,.Q6(Q[1517])			,.R1(R[1512])	,.R2(R[1513])	,.R3(R[1514])	,.R4(R[1515])	,.R5(R[1516])	,.R6(R[1517])			,.clk(clk)	);
CNU_6 CNU238	(.Q1(Q[1518])	,.Q2(Q[1519])	,.Q3(Q[1520])	,.Q4(Q[1521])	,.Q5(Q[1522])	,.Q6(Q[1523])			,.R1(R[1518])	,.R2(R[1519])	,.R3(R[1520])	,.R4(R[1521])	,.R5(R[1522])	,.R6(R[1523])			,.clk(clk)	);
CNU_6 CNU239	(.Q1(Q[1524])	,.Q2(Q[1525])	,.Q3(Q[1526])	,.Q4(Q[1527])	,.Q5(Q[1528])	,.Q6(Q[1529])			,.R1(R[1524])	,.R2(R[1525])	,.R3(R[1526])	,.R4(R[1527])	,.R5(R[1528])	,.R6(R[1529])			,.clk(clk)	);
CNU_6 CNU240	(.Q1(Q[1530])	,.Q2(Q[1531])	,.Q3(Q[1532])	,.Q4(Q[1533])	,.Q5(Q[1534])	,.Q6(Q[1535])			,.R1(R[1530])	,.R2(R[1531])	,.R3(R[1532])	,.R4(R[1533])	,.R5(R[1534])	,.R6(R[1535])			,.clk(clk)	);
CNU_6 CNU241	(.Q1(Q[1536])	,.Q2(Q[1537])	,.Q3(Q[1538])	,.Q4(Q[1539])	,.Q5(Q[1540])	,.Q6(Q[1541])			,.R1(R[1536])	,.R2(R[1537])	,.R3(R[1538])	,.R4(R[1539])	,.R5(R[1540])	,.R6(R[1541])			,.clk(clk)	);
CNU_6 CNU242	(.Q1(Q[1542])	,.Q2(Q[1543])	,.Q3(Q[1544])	,.Q4(Q[1545])	,.Q5(Q[1546])	,.Q6(Q[1547])			,.R1(R[1542])	,.R2(R[1543])	,.R3(R[1544])	,.R4(R[1545])	,.R5(R[1546])	,.R6(R[1547])			,.clk(clk)	);
CNU_6 CNU243	(.Q1(Q[1548])	,.Q2(Q[1549])	,.Q3(Q[1550])	,.Q4(Q[1551])	,.Q5(Q[1552])	,.Q6(Q[1553])			,.R1(R[1548])	,.R2(R[1549])	,.R3(R[1550])	,.R4(R[1551])	,.R5(R[1552])	,.R6(R[1553])			,.clk(clk)	);
CNU_6 CNU244	(.Q1(Q[1554])	,.Q2(Q[1555])	,.Q3(Q[1556])	,.Q4(Q[1557])	,.Q5(Q[1558])	,.Q6(Q[1559])			,.R1(R[1554])	,.R2(R[1555])	,.R3(R[1556])	,.R4(R[1557])	,.R5(R[1558])	,.R6(R[1559])			,.clk(clk)	);
CNU_6 CNU245	(.Q1(Q[1560])	,.Q2(Q[1561])	,.Q3(Q[1562])	,.Q4(Q[1563])	,.Q5(Q[1564])	,.Q6(Q[1565])			,.R1(R[1560])	,.R2(R[1561])	,.R3(R[1562])	,.R4(R[1563])	,.R5(R[1564])	,.R6(R[1565])			,.clk(clk)	);
CNU_6 CNU246	(.Q1(Q[1566])	,.Q2(Q[1567])	,.Q3(Q[1568])	,.Q4(Q[1569])	,.Q5(Q[1570])	,.Q6(Q[1571])			,.R1(R[1566])	,.R2(R[1567])	,.R3(R[1568])	,.R4(R[1569])	,.R5(R[1570])	,.R6(R[1571])			,.clk(clk)	);
CNU_6 CNU247	(.Q1(Q[1572])	,.Q2(Q[1573])	,.Q3(Q[1574])	,.Q4(Q[1575])	,.Q5(Q[1576])	,.Q6(Q[1577])			,.R1(R[1572])	,.R2(R[1573])	,.R3(R[1574])	,.R4(R[1575])	,.R5(R[1576])	,.R6(R[1577])			,.clk(clk)	);
CNU_6 CNU248	(.Q1(Q[1578])	,.Q2(Q[1579])	,.Q3(Q[1580])	,.Q4(Q[1581])	,.Q5(Q[1582])	,.Q6(Q[1583])			,.R1(R[1578])	,.R2(R[1579])	,.R3(R[1580])	,.R4(R[1581])	,.R5(R[1582])	,.R6(R[1583])			,.clk(clk)	);
CNU_6 CNU249	(.Q1(Q[1584])	,.Q2(Q[1585])	,.Q3(Q[1586])	,.Q4(Q[1587])	,.Q5(Q[1588])	,.Q6(Q[1589])			,.R1(R[1584])	,.R2(R[1585])	,.R3(R[1586])	,.R4(R[1587])	,.R5(R[1588])	,.R6(R[1589])			,.clk(clk)	);
CNU_6 CNU250	(.Q1(Q[1590])	,.Q2(Q[1591])	,.Q3(Q[1592])	,.Q4(Q[1593])	,.Q5(Q[1594])	,.Q6(Q[1595])			,.R1(R[1590])	,.R2(R[1591])	,.R3(R[1592])	,.R4(R[1593])	,.R5(R[1594])	,.R6(R[1595])			,.clk(clk)	);
CNU_6 CNU251	(.Q1(Q[1596])	,.Q2(Q[1597])	,.Q3(Q[1598])	,.Q4(Q[1599])	,.Q5(Q[1600])	,.Q6(Q[1601])			,.R1(R[1596])	,.R2(R[1597])	,.R3(R[1598])	,.R4(R[1599])	,.R5(R[1600])	,.R6(R[1601])			,.clk(clk)	);
CNU_6 CNU252	(.Q1(Q[1602])	,.Q2(Q[1603])	,.Q3(Q[1604])	,.Q4(Q[1605])	,.Q5(Q[1606])	,.Q6(Q[1607])			,.R1(R[1602])	,.R2(R[1603])	,.R3(R[1604])	,.R4(R[1605])	,.R5(R[1606])	,.R6(R[1607])			,.clk(clk)	);
CNU_6 CNU253	(.Q1(Q[1608])	,.Q2(Q[1609])	,.Q3(Q[1610])	,.Q4(Q[1611])	,.Q5(Q[1612])	,.Q6(Q[1613])			,.R1(R[1608])	,.R2(R[1609])	,.R3(R[1610])	,.R4(R[1611])	,.R5(R[1612])	,.R6(R[1613])			,.clk(clk)	);
CNU_6 CNU254	(.Q1(Q[1614])	,.Q2(Q[1615])	,.Q3(Q[1616])	,.Q4(Q[1617])	,.Q5(Q[1618])	,.Q6(Q[1619])			,.R1(R[1614])	,.R2(R[1615])	,.R3(R[1616])	,.R4(R[1617])	,.R5(R[1618])	,.R6(R[1619])			,.clk(clk)	);
CNU_6 CNU255	(.Q1(Q[1620])	,.Q2(Q[1621])	,.Q3(Q[1622])	,.Q4(Q[1623])	,.Q5(Q[1624])	,.Q6(Q[1625])			,.R1(R[1620])	,.R2(R[1621])	,.R3(R[1622])	,.R4(R[1623])	,.R5(R[1624])	,.R6(R[1625])			,.clk(clk)	);
CNU_6 CNU256	(.Q1(Q[1626])	,.Q2(Q[1627])	,.Q3(Q[1628])	,.Q4(Q[1629])	,.Q5(Q[1630])	,.Q6(Q[1631])			,.R1(R[1626])	,.R2(R[1627])	,.R3(R[1628])	,.R4(R[1629])	,.R5(R[1630])	,.R6(R[1631])			,.clk(clk)	);
CNU_6 CNU257	(.Q1(Q[1632])	,.Q2(Q[1633])	,.Q3(Q[1634])	,.Q4(Q[1635])	,.Q5(Q[1636])	,.Q6(Q[1637])			,.R1(R[1632])	,.R2(R[1633])	,.R3(R[1634])	,.R4(R[1635])	,.R5(R[1636])	,.R6(R[1637])			,.clk(clk)	);
CNU_6 CNU258	(.Q1(Q[1638])	,.Q2(Q[1639])	,.Q3(Q[1640])	,.Q4(Q[1641])	,.Q5(Q[1642])	,.Q6(Q[1643])			,.R1(R[1638])	,.R2(R[1639])	,.R3(R[1640])	,.R4(R[1641])	,.R5(R[1642])	,.R6(R[1643])			,.clk(clk)	);
CNU_6 CNU259	(.Q1(Q[1644])	,.Q2(Q[1645])	,.Q3(Q[1646])	,.Q4(Q[1647])	,.Q5(Q[1648])	,.Q6(Q[1649])			,.R1(R[1644])	,.R2(R[1645])	,.R3(R[1646])	,.R4(R[1647])	,.R5(R[1648])	,.R6(R[1649])			,.clk(clk)	);
CNU_6 CNU260	(.Q1(Q[1650])	,.Q2(Q[1651])	,.Q3(Q[1652])	,.Q4(Q[1653])	,.Q5(Q[1654])	,.Q6(Q[1655])			,.R1(R[1650])	,.R2(R[1651])	,.R3(R[1652])	,.R4(R[1653])	,.R5(R[1654])	,.R6(R[1655])			,.clk(clk)	);
CNU_6 CNU261	(.Q1(Q[1656])	,.Q2(Q[1657])	,.Q3(Q[1658])	,.Q4(Q[1659])	,.Q5(Q[1660])	,.Q6(Q[1661])			,.R1(R[1656])	,.R2(R[1657])	,.R3(R[1658])	,.R4(R[1659])	,.R5(R[1660])	,.R6(R[1661])			,.clk(clk)	);
CNU_6 CNU262	(.Q1(Q[1662])	,.Q2(Q[1663])	,.Q3(Q[1664])	,.Q4(Q[1665])	,.Q5(Q[1666])	,.Q6(Q[1667])			,.R1(R[1662])	,.R2(R[1663])	,.R3(R[1664])	,.R4(R[1665])	,.R5(R[1666])	,.R6(R[1667])			,.clk(clk)	);
CNU_6 CNU263	(.Q1(Q[1668])	,.Q2(Q[1669])	,.Q3(Q[1670])	,.Q4(Q[1671])	,.Q5(Q[1672])	,.Q6(Q[1673])			,.R1(R[1668])	,.R2(R[1669])	,.R3(R[1670])	,.R4(R[1671])	,.R5(R[1672])	,.R6(R[1673])			,.clk(clk)	);
CNU_6 CNU264	(.Q1(Q[1674])	,.Q2(Q[1675])	,.Q3(Q[1676])	,.Q4(Q[1677])	,.Q5(Q[1678])	,.Q6(Q[1679])			,.R1(R[1674])	,.R2(R[1675])	,.R3(R[1676])	,.R4(R[1677])	,.R5(R[1678])	,.R6(R[1679])			,.clk(clk)	);
CNU_6 CNU265	(.Q1(Q[1680])	,.Q2(Q[1681])	,.Q3(Q[1682])	,.Q4(Q[1683])	,.Q5(Q[1684])	,.Q6(Q[1685])			,.R1(R[1680])	,.R2(R[1681])	,.R3(R[1682])	,.R4(R[1683])	,.R5(R[1684])	,.R6(R[1685])			,.clk(clk)	);
CNU_6 CNU266	(.Q1(Q[1686])	,.Q2(Q[1687])	,.Q3(Q[1688])	,.Q4(Q[1689])	,.Q5(Q[1690])	,.Q6(Q[1691])			,.R1(R[1686])	,.R2(R[1687])	,.R3(R[1688])	,.R4(R[1689])	,.R5(R[1690])	,.R6(R[1691])			,.clk(clk)	);
CNU_6 CNU267	(.Q1(Q[1692])	,.Q2(Q[1693])	,.Q3(Q[1694])	,.Q4(Q[1695])	,.Q5(Q[1696])	,.Q6(Q[1697])			,.R1(R[1692])	,.R2(R[1693])	,.R3(R[1694])	,.R4(R[1695])	,.R5(R[1696])	,.R6(R[1697])			,.clk(clk)	);
CNU_6 CNU268	(.Q1(Q[1698])	,.Q2(Q[1699])	,.Q3(Q[1700])	,.Q4(Q[1701])	,.Q5(Q[1702])	,.Q6(Q[1703])			,.R1(R[1698])	,.R2(R[1699])	,.R3(R[1700])	,.R4(R[1701])	,.R5(R[1702])	,.R6(R[1703])			,.clk(clk)	);
CNU_6 CNU269	(.Q1(Q[1704])	,.Q2(Q[1705])	,.Q3(Q[1706])	,.Q4(Q[1707])	,.Q5(Q[1708])	,.Q6(Q[1709])			,.R1(R[1704])	,.R2(R[1705])	,.R3(R[1706])	,.R4(R[1707])	,.R5(R[1708])	,.R6(R[1709])			,.clk(clk)	);
CNU_6 CNU270	(.Q1(Q[1710])	,.Q2(Q[1711])	,.Q3(Q[1712])	,.Q4(Q[1713])	,.Q5(Q[1714])	,.Q6(Q[1715])			,.R1(R[1710])	,.R2(R[1711])	,.R3(R[1712])	,.R4(R[1713])	,.R5(R[1714])	,.R6(R[1715])			,.clk(clk)	);
CNU_6 CNU271	(.Q1(Q[1716])	,.Q2(Q[1717])	,.Q3(Q[1718])	,.Q4(Q[1719])	,.Q5(Q[1720])	,.Q6(Q[1721])			,.R1(R[1716])	,.R2(R[1717])	,.R3(R[1718])	,.R4(R[1719])	,.R5(R[1720])	,.R6(R[1721])			,.clk(clk)	);
CNU_6 CNU272	(.Q1(Q[1722])	,.Q2(Q[1723])	,.Q3(Q[1724])	,.Q4(Q[1725])	,.Q5(Q[1726])	,.Q6(Q[1727])			,.R1(R[1722])	,.R2(R[1723])	,.R3(R[1724])	,.R4(R[1725])	,.R5(R[1726])	,.R6(R[1727])			,.clk(clk)	);
CNU_6 CNU273	(.Q1(Q[1728])	,.Q2(Q[1729])	,.Q3(Q[1730])	,.Q4(Q[1731])	,.Q5(Q[1732])	,.Q6(Q[1733])			,.R1(R[1728])	,.R2(R[1729])	,.R3(R[1730])	,.R4(R[1731])	,.R5(R[1732])	,.R6(R[1733])			,.clk(clk)	);
CNU_6 CNU274	(.Q1(Q[1734])	,.Q2(Q[1735])	,.Q3(Q[1736])	,.Q4(Q[1737])	,.Q5(Q[1738])	,.Q6(Q[1739])			,.R1(R[1734])	,.R2(R[1735])	,.R3(R[1736])	,.R4(R[1737])	,.R5(R[1738])	,.R6(R[1739])			,.clk(clk)	);
CNU_6 CNU275	(.Q1(Q[1740])	,.Q2(Q[1741])	,.Q3(Q[1742])	,.Q4(Q[1743])	,.Q5(Q[1744])	,.Q6(Q[1745])			,.R1(R[1740])	,.R2(R[1741])	,.R3(R[1742])	,.R4(R[1743])	,.R5(R[1744])	,.R6(R[1745])			,.clk(clk)	);
CNU_6 CNU276	(.Q1(Q[1746])	,.Q2(Q[1747])	,.Q3(Q[1748])	,.Q4(Q[1749])	,.Q5(Q[1750])	,.Q6(Q[1751])			,.R1(R[1746])	,.R2(R[1747])	,.R3(R[1748])	,.R4(R[1749])	,.R5(R[1750])	,.R6(R[1751])			,.clk(clk)	);
CNU_6 CNU277	(.Q1(Q[1752])	,.Q2(Q[1753])	,.Q3(Q[1754])	,.Q4(Q[1755])	,.Q5(Q[1756])	,.Q6(Q[1757])			,.R1(R[1752])	,.R2(R[1753])	,.R3(R[1754])	,.R4(R[1755])	,.R5(R[1756])	,.R6(R[1757])			,.clk(clk)	);
CNU_6 CNU278	(.Q1(Q[1758])	,.Q2(Q[1759])	,.Q3(Q[1760])	,.Q4(Q[1761])	,.Q5(Q[1762])	,.Q6(Q[1763])			,.R1(R[1758])	,.R2(R[1759])	,.R3(R[1760])	,.R4(R[1761])	,.R5(R[1762])	,.R6(R[1763])			,.clk(clk)	);
CNU_6 CNU279	(.Q1(Q[1764])	,.Q2(Q[1765])	,.Q3(Q[1766])	,.Q4(Q[1767])	,.Q5(Q[1768])	,.Q6(Q[1769])			,.R1(R[1764])	,.R2(R[1765])	,.R3(R[1766])	,.R4(R[1767])	,.R5(R[1768])	,.R6(R[1769])			,.clk(clk)	);
CNU_6 CNU280	(.Q1(Q[1770])	,.Q2(Q[1771])	,.Q3(Q[1772])	,.Q4(Q[1773])	,.Q5(Q[1774])	,.Q6(Q[1775])			,.R1(R[1770])	,.R2(R[1771])	,.R3(R[1772])	,.R4(R[1773])	,.R5(R[1774])	,.R6(R[1775])			,.clk(clk)	);
CNU_6 CNU281	(.Q1(Q[1776])	,.Q2(Q[1777])	,.Q3(Q[1778])	,.Q4(Q[1779])	,.Q5(Q[1780])	,.Q6(Q[1781])			,.R1(R[1776])	,.R2(R[1777])	,.R3(R[1778])	,.R4(R[1779])	,.R5(R[1780])	,.R6(R[1781])			,.clk(clk)	);
CNU_6 CNU282	(.Q1(Q[1782])	,.Q2(Q[1783])	,.Q3(Q[1784])	,.Q4(Q[1785])	,.Q5(Q[1786])	,.Q6(Q[1787])			,.R1(R[1782])	,.R2(R[1783])	,.R3(R[1784])	,.R4(R[1785])	,.R5(R[1786])	,.R6(R[1787])			,.clk(clk)	);
CNU_6 CNU283	(.Q1(Q[1788])	,.Q2(Q[1789])	,.Q3(Q[1790])	,.Q4(Q[1791])	,.Q5(Q[1792])	,.Q6(Q[1793])			,.R1(R[1788])	,.R2(R[1789])	,.R3(R[1790])	,.R4(R[1791])	,.R5(R[1792])	,.R6(R[1793])			,.clk(clk)	);
CNU_6 CNU284	(.Q1(Q[1794])	,.Q2(Q[1795])	,.Q3(Q[1796])	,.Q4(Q[1797])	,.Q5(Q[1798])	,.Q6(Q[1799])			,.R1(R[1794])	,.R2(R[1795])	,.R3(R[1796])	,.R4(R[1797])	,.R5(R[1798])	,.R6(R[1799])			,.clk(clk)	);
CNU_6 CNU285	(.Q1(Q[1800])	,.Q2(Q[1801])	,.Q3(Q[1802])	,.Q4(Q[1803])	,.Q5(Q[1804])	,.Q6(Q[1805])			,.R1(R[1800])	,.R2(R[1801])	,.R3(R[1802])	,.R4(R[1803])	,.R5(R[1804])	,.R6(R[1805])			,.clk(clk)	);
CNU_6 CNU286	(.Q1(Q[1806])	,.Q2(Q[1807])	,.Q3(Q[1808])	,.Q4(Q[1809])	,.Q5(Q[1810])	,.Q6(Q[1811])			,.R1(R[1806])	,.R2(R[1807])	,.R3(R[1808])	,.R4(R[1809])	,.R5(R[1810])	,.R6(R[1811])			,.clk(clk)	);
CNU_6 CNU287	(.Q1(Q[1812])	,.Q2(Q[1813])	,.Q3(Q[1814])	,.Q4(Q[1815])	,.Q5(Q[1816])	,.Q6(Q[1817])			,.R1(R[1812])	,.R2(R[1813])	,.R3(R[1814])	,.R4(R[1815])	,.R5(R[1816])	,.R6(R[1817])			,.clk(clk)	);
CNU_6 CNU288	(.Q1(Q[1818])	,.Q2(Q[1819])	,.Q3(Q[1820])	,.Q4(Q[1821])	,.Q5(Q[1822])	,.Q6(Q[1823])			,.R1(R[1818])	,.R2(R[1819])	,.R3(R[1820])	,.R4(R[1821])	,.R5(R[1822])	,.R6(R[1823])			,.clk(clk)	);


VNU_3 VNU1	(.Q1(Q[534])	,.Q2(Q[1371])	,.Q3(Q[1764])							,.R1(R[534])	,.R2(R[1371])	,.R3(R[1764])							,.clk(clk)	,.L(L1)	,.P(P[0])	,.reset(reset)	);
VNU_3 VNU2	(.Q1(Q[540])	,.Q2(Q[1378])	,.Q3(Q[1770])							,.R1(R[540])	,.R2(R[1378])	,.R3(R[1770])							,.clk(clk)	,.L(L2)	,.P(P[1])	,.reset(reset)	);
VNU_3 VNU3	(.Q1(Q[546])	,.Q2(Q[1385])	,.Q3(Q[1776])							,.R1(R[546])	,.R2(R[1385])	,.R3(R[1776])							,.clk(clk)	,.L(L3)	,.P(P[2])	,.reset(reset)	);
VNU_3 VNU4	(.Q1(Q[552])	,.Q2(Q[1224])	,.Q3(Q[1782])							,.R1(R[552])	,.R2(R[1224])	,.R3(R[1782])							,.clk(clk)	,.L(L4)	,.P(P[3])	,.reset(reset)	);
VNU_3 VNU5	(.Q1(Q[558])	,.Q2(Q[1231])	,.Q3(Q[1788])							,.R1(R[558])	,.R2(R[1231])	,.R3(R[1788])							,.clk(clk)	,.L(L5)	,.P(P[4])	,.reset(reset)	);
VNU_3 VNU6	(.Q1(Q[564])	,.Q2(Q[1238])	,.Q3(Q[1794])							,.R1(R[564])	,.R2(R[1238])	,.R3(R[1794])							,.clk(clk)	,.L(L6)	,.P(P[5])	,.reset(reset)	);
VNU_3 VNU7	(.Q1(Q[570])	,.Q2(Q[1245])	,.Q3(Q[1800])							,.R1(R[570])	,.R2(R[1245])	,.R3(R[1800])							,.clk(clk)	,.L(L7)	,.P(P[6])	,.reset(reset)	);
VNU_3 VNU8	(.Q1(Q[576])	,.Q2(Q[1252])	,.Q3(Q[1806])							,.R1(R[576])	,.R2(R[1252])	,.R3(R[1806])							,.clk(clk)	,.L(L8)	,.P(P[7])	,.reset(reset)	);
VNU_3 VNU9	(.Q1(Q[582])	,.Q2(Q[1259])	,.Q3(Q[1812])							,.R1(R[582])	,.R2(R[1259])	,.R3(R[1812])							,.clk(clk)	,.L(L9)	,.P(P[8])	,.reset(reset)	);
VNU_3 VNU10	(.Q1(Q[588])	,.Q2(Q[1266])	,.Q3(Q[1818])							,.R1(R[588])	,.R2(R[1266])	,.R3(R[1818])							,.clk(clk)	,.L(L10)	,.P(P[9])	,.reset(reset)	);
VNU_3 VNU11	(.Q1(Q[594])	,.Q2(Q[1273])	,.Q3(Q[1680])							,.R1(R[594])	,.R2(R[1273])	,.R3(R[1680])							,.clk(clk)	,.L(L11)	,.P(P[10])	,.reset(reset)	);
VNU_3 VNU12	(.Q1(Q[600])	,.Q2(Q[1280])	,.Q3(Q[1686])							,.R1(R[600])	,.R2(R[1280])	,.R3(R[1686])							,.clk(clk)	,.L(L12)	,.P(P[11])	,.reset(reset)	);
VNU_3 VNU13	(.Q1(Q[606])	,.Q2(Q[1287])	,.Q3(Q[1692])							,.R1(R[606])	,.R2(R[1287])	,.R3(R[1692])							,.clk(clk)	,.L(L13)	,.P(P[12])	,.reset(reset)	);
VNU_3 VNU14	(.Q1(Q[612])	,.Q2(Q[1294])	,.Q3(Q[1698])							,.R1(R[612])	,.R2(R[1294])	,.R3(R[1698])							,.clk(clk)	,.L(L14)	,.P(P[13])	,.reset(reset)	);
VNU_3 VNU15	(.Q1(Q[618])	,.Q2(Q[1301])	,.Q3(Q[1704])							,.R1(R[618])	,.R2(R[1301])	,.R3(R[1704])							,.clk(clk)	,.L(L15)	,.P(P[14])	,.reset(reset)	);
VNU_3 VNU16	(.Q1(Q[480])	,.Q2(Q[1308])	,.Q3(Q[1710])							,.R1(R[480])	,.R2(R[1308])	,.R3(R[1710])							,.clk(clk)	,.L(L16)	,.P(P[15])	,.reset(reset)	);
VNU_3 VNU17	(.Q1(Q[486])	,.Q2(Q[1315])	,.Q3(Q[1716])							,.R1(R[486])	,.R2(R[1315])	,.R3(R[1716])							,.clk(clk)	,.L(L17)	,.P(P[16])	,.reset(reset)	);
VNU_3 VNU18	(.Q1(Q[492])	,.Q2(Q[1322])	,.Q3(Q[1722])							,.R1(R[492])	,.R2(R[1322])	,.R3(R[1722])							,.clk(clk)	,.L(L18)	,.P(P[17])	,.reset(reset)	);
VNU_3 VNU19	(.Q1(Q[498])	,.Q2(Q[1329])	,.Q3(Q[1728])							,.R1(R[498])	,.R2(R[1329])	,.R3(R[1728])							,.clk(clk)	,.L(L19)	,.P(P[18])	,.reset(reset)	);
VNU_3 VNU20	(.Q1(Q[504])	,.Q2(Q[1336])	,.Q3(Q[1734])							,.R1(R[504])	,.R2(R[1336])	,.R3(R[1734])							,.clk(clk)	,.L(L20)	,.P(P[19])	,.reset(reset)	);
VNU_3 VNU21	(.Q1(Q[510])	,.Q2(Q[1343])	,.Q3(Q[1740])							,.R1(R[510])	,.R2(R[1343])	,.R3(R[1740])							,.clk(clk)	,.L(L21)	,.P(P[20])	,.reset(reset)	);
VNU_3 VNU22	(.Q1(Q[516])	,.Q2(Q[1350])	,.Q3(Q[1746])							,.R1(R[516])	,.R2(R[1350])	,.R3(R[1746])							,.clk(clk)	,.L(L22)	,.P(P[21])	,.reset(reset)	);
VNU_3 VNU23	(.Q1(Q[522])	,.Q2(Q[1357])	,.Q3(Q[1752])							,.R1(R[522])	,.R2(R[1357])	,.R3(R[1752])							,.clk(clk)	,.L(L23)	,.P(P[22])	,.reset(reset)	);
VNU_3 VNU24	(.Q1(Q[528])	,.Q2(Q[1364])	,.Q3(Q[1758])							,.R1(R[528])	,.R2(R[1364])	,.R3(R[1758])							,.clk(clk)	,.L(L24)	,.P(P[23])	,.reset(reset)	);
VNU_3 VNU25	(.Q1(Q[6])	,.Q2(Q[270])	,.Q3(Q[1212])							,.R1(R[6])	,.R2(R[270])	,.R3(R[1212])							,.clk(clk)	,.L(L25)	,.P(P[24])	,.reset(reset)	);
VNU_3 VNU26	(.Q1(Q[12])	,.Q2(Q[277])	,.Q3(Q[1218])							,.R1(R[12])	,.R2(R[277])	,.R3(R[1218])							,.clk(clk)	,.L(L26)	,.P(P[25])	,.reset(reset)	);
VNU_3 VNU27	(.Q1(Q[18])	,.Q2(Q[284])	,.Q3(Q[1080])							,.R1(R[18])	,.R2(R[284])	,.R3(R[1080])							,.clk(clk)	,.L(L27)	,.P(P[26])	,.reset(reset)	);
VNU_3 VNU28	(.Q1(Q[24])	,.Q2(Q[291])	,.Q3(Q[1086])							,.R1(R[24])	,.R2(R[291])	,.R3(R[1086])							,.clk(clk)	,.L(L28)	,.P(P[27])	,.reset(reset)	);
VNU_3 VNU29	(.Q1(Q[30])	,.Q2(Q[298])	,.Q3(Q[1092])							,.R1(R[30])	,.R2(R[298])	,.R3(R[1092])							,.clk(clk)	,.L(L29)	,.P(P[28])	,.reset(reset)	);
VNU_3 VNU30	(.Q1(Q[36])	,.Q2(Q[305])	,.Q3(Q[1098])							,.R1(R[36])	,.R2(R[305])	,.R3(R[1098])							,.clk(clk)	,.L(L30)	,.P(P[29])	,.reset(reset)	);
VNU_3 VNU31	(.Q1(Q[42])	,.Q2(Q[144])	,.Q3(Q[1104])							,.R1(R[42])	,.R2(R[144])	,.R3(R[1104])							,.clk(clk)	,.L(L31)	,.P(P[30])	,.reset(reset)	);
VNU_3 VNU32	(.Q1(Q[48])	,.Q2(Q[151])	,.Q3(Q[1110])							,.R1(R[48])	,.R2(R[151])	,.R3(R[1110])							,.clk(clk)	,.L(L32)	,.P(P[31])	,.reset(reset)	);
VNU_3 VNU33	(.Q1(Q[54])	,.Q2(Q[158])	,.Q3(Q[1116])							,.R1(R[54])	,.R2(R[158])	,.R3(R[1116])							,.clk(clk)	,.L(L33)	,.P(P[32])	,.reset(reset)	);
VNU_3 VNU34	(.Q1(Q[60])	,.Q2(Q[165])	,.Q3(Q[1122])							,.R1(R[60])	,.R2(R[165])	,.R3(R[1122])							,.clk(clk)	,.L(L34)	,.P(P[33])	,.reset(reset)	);
VNU_3 VNU35	(.Q1(Q[66])	,.Q2(Q[172])	,.Q3(Q[1128])							,.R1(R[66])	,.R2(R[172])	,.R3(R[1128])							,.clk(clk)	,.L(L35)	,.P(P[34])	,.reset(reset)	);
VNU_3 VNU36	(.Q1(Q[72])	,.Q2(Q[179])	,.Q3(Q[1134])							,.R1(R[72])	,.R2(R[179])	,.R3(R[1134])							,.clk(clk)	,.L(L36)	,.P(P[35])	,.reset(reset)	);
VNU_3 VNU37	(.Q1(Q[78])	,.Q2(Q[186])	,.Q3(Q[1140])							,.R1(R[78])	,.R2(R[186])	,.R3(R[1140])							,.clk(clk)	,.L(L37)	,.P(P[36])	,.reset(reset)	);
VNU_3 VNU38	(.Q1(Q[84])	,.Q2(Q[193])	,.Q3(Q[1146])							,.R1(R[84])	,.R2(R[193])	,.R3(R[1146])							,.clk(clk)	,.L(L38)	,.P(P[37])	,.reset(reset)	);
VNU_3 VNU39	(.Q1(Q[90])	,.Q2(Q[200])	,.Q3(Q[1152])							,.R1(R[90])	,.R2(R[200])	,.R3(R[1152])							,.clk(clk)	,.L(L39)	,.P(P[38])	,.reset(reset)	);
VNU_3 VNU40	(.Q1(Q[96])	,.Q2(Q[207])	,.Q3(Q[1158])							,.R1(R[96])	,.R2(R[207])	,.R3(R[1158])							,.clk(clk)	,.L(L40)	,.P(P[39])	,.reset(reset)	);
VNU_3 VNU41	(.Q1(Q[102])	,.Q2(Q[214])	,.Q3(Q[1164])							,.R1(R[102])	,.R2(R[214])	,.R3(R[1164])							,.clk(clk)	,.L(L41)	,.P(P[40])	,.reset(reset)	);
VNU_3 VNU42	(.Q1(Q[108])	,.Q2(Q[221])	,.Q3(Q[1170])							,.R1(R[108])	,.R2(R[221])	,.R3(R[1170])							,.clk(clk)	,.L(L42)	,.P(P[41])	,.reset(reset)	);
VNU_3 VNU43	(.Q1(Q[114])	,.Q2(Q[228])	,.Q3(Q[1176])							,.R1(R[114])	,.R2(R[228])	,.R3(R[1176])							,.clk(clk)	,.L(L43)	,.P(P[42])	,.reset(reset)	);
VNU_3 VNU44	(.Q1(Q[120])	,.Q2(Q[235])	,.Q3(Q[1182])							,.R1(R[120])	,.R2(R[235])	,.R3(R[1182])							,.clk(clk)	,.L(L44)	,.P(P[43])	,.reset(reset)	);
VNU_3 VNU45	(.Q1(Q[126])	,.Q2(Q[242])	,.Q3(Q[1188])							,.R1(R[126])	,.R2(R[242])	,.R3(R[1188])							,.clk(clk)	,.L(L45)	,.P(P[44])	,.reset(reset)	);
VNU_3 VNU46	(.Q1(Q[132])	,.Q2(Q[249])	,.Q3(Q[1194])							,.R1(R[132])	,.R2(R[249])	,.R3(R[1194])							,.clk(clk)	,.L(L46)	,.P(P[45])	,.reset(reset)	);
VNU_3 VNU47	(.Q1(Q[138])	,.Q2(Q[256])	,.Q3(Q[1200])							,.R1(R[138])	,.R2(R[256])	,.R3(R[1200])							,.clk(clk)	,.L(L47)	,.P(P[46])	,.reset(reset)	);
VNU_3 VNU48	(.Q1(Q[0])	,.Q2(Q[263])	,.Q3(Q[1206])							,.R1(R[0])	,.R2(R[263])	,.R3(R[1206])							,.clk(clk)	,.L(L48)	,.P(P[47])	,.reset(reset)	);
VNU_6 VNU49	(.Q1(Q[37])	,.Q2(Q[559])	,.Q3(Q[714])	,.Q4(Q[942])	,.Q5(Q[1117])	,.Q6(Q[1674])	,.R1(R[37])	,.R2(R[559])	,.R3(R[714])	,.R4(R[942])	,.R5(R[1117])	,.R6(R[1674])	,.clk(clk)	,.L(L49)	,.P(P[48])	,.reset(reset)	);
VNU_6 VNU50	(.Q1(Q[43])	,.Q2(Q[565])	,.Q3(Q[720])	,.Q4(Q[948])	,.Q5(Q[1123])	,.Q6(Q[1536])	,.R1(R[43])	,.R2(R[565])	,.R3(R[720])	,.R4(R[948])	,.R5(R[1123])	,.R6(R[1536])	,.clk(clk)	,.L(L50)	,.P(P[49])	,.reset(reset)	);
VNU_6 VNU51	(.Q1(Q[49])	,.Q2(Q[571])	,.Q3(Q[726])	,.Q4(Q[954])	,.Q5(Q[1129])	,.Q6(Q[1542])	,.R1(R[49])	,.R2(R[571])	,.R3(R[726])	,.R4(R[954])	,.R5(R[1129])	,.R6(R[1542])	,.clk(clk)	,.L(L51)	,.P(P[50])	,.reset(reset)	);
VNU_6 VNU52	(.Q1(Q[55])	,.Q2(Q[577])	,.Q3(Q[732])	,.Q4(Q[960])	,.Q5(Q[1135])	,.Q6(Q[1548])	,.R1(R[55])	,.R2(R[577])	,.R3(R[732])	,.R4(R[960])	,.R5(R[1135])	,.R6(R[1548])	,.clk(clk)	,.L(L52)	,.P(P[51])	,.reset(reset)	);
VNU_6 VNU53	(.Q1(Q[61])	,.Q2(Q[583])	,.Q3(Q[738])	,.Q4(Q[966])	,.Q5(Q[1141])	,.Q6(Q[1554])	,.R1(R[61])	,.R2(R[583])	,.R3(R[738])	,.R4(R[966])	,.R5(R[1141])	,.R6(R[1554])	,.clk(clk)	,.L(L53)	,.P(P[52])	,.reset(reset)	);
VNU_6 VNU54	(.Q1(Q[67])	,.Q2(Q[589])	,.Q3(Q[744])	,.Q4(Q[972])	,.Q5(Q[1147])	,.Q6(Q[1560])	,.R1(R[67])	,.R2(R[589])	,.R3(R[744])	,.R4(R[972])	,.R5(R[1147])	,.R6(R[1560])	,.clk(clk)	,.L(L54)	,.P(P[53])	,.reset(reset)	);
VNU_6 VNU55	(.Q1(Q[73])	,.Q2(Q[595])	,.Q3(Q[750])	,.Q4(Q[978])	,.Q5(Q[1153])	,.Q6(Q[1566])	,.R1(R[73])	,.R2(R[595])	,.R3(R[750])	,.R4(R[978])	,.R5(R[1153])	,.R6(R[1566])	,.clk(clk)	,.L(L55)	,.P(P[54])	,.reset(reset)	);
VNU_6 VNU56	(.Q1(Q[79])	,.Q2(Q[601])	,.Q3(Q[756])	,.Q4(Q[984])	,.Q5(Q[1159])	,.Q6(Q[1572])	,.R1(R[79])	,.R2(R[601])	,.R3(R[756])	,.R4(R[984])	,.R5(R[1159])	,.R6(R[1572])	,.clk(clk)	,.L(L56)	,.P(P[55])	,.reset(reset)	);
VNU_6 VNU57	(.Q1(Q[85])	,.Q2(Q[607])	,.Q3(Q[762])	,.Q4(Q[990])	,.Q5(Q[1165])	,.Q6(Q[1578])	,.R1(R[85])	,.R2(R[607])	,.R3(R[762])	,.R4(R[990])	,.R5(R[1165])	,.R6(R[1578])	,.clk(clk)	,.L(L57)	,.P(P[56])	,.reset(reset)	);
VNU_6 VNU58	(.Q1(Q[91])	,.Q2(Q[613])	,.Q3(Q[624])	,.Q4(Q[996])	,.Q5(Q[1171])	,.Q6(Q[1584])	,.R1(R[91])	,.R2(R[613])	,.R3(R[624])	,.R4(R[996])	,.R5(R[1171])	,.R6(R[1584])	,.clk(clk)	,.L(L58)	,.P(P[57])	,.reset(reset)	);
VNU_6 VNU59	(.Q1(Q[97])	,.Q2(Q[619])	,.Q3(Q[630])	,.Q4(Q[1002])	,.Q5(Q[1177])	,.Q6(Q[1590])	,.R1(R[97])	,.R2(R[619])	,.R3(R[630])	,.R4(R[1002])	,.R5(R[1177])	,.R6(R[1590])	,.clk(clk)	,.L(L59)	,.P(P[58])	,.reset(reset)	);
VNU_6 VNU60	(.Q1(Q[103])	,.Q2(Q[481])	,.Q3(Q[636])	,.Q4(Q[1008])	,.Q5(Q[1183])	,.Q6(Q[1596])	,.R1(R[103])	,.R2(R[481])	,.R3(R[636])	,.R4(R[1008])	,.R5(R[1183])	,.R6(R[1596])	,.clk(clk)	,.L(L60)	,.P(P[59])	,.reset(reset)	);
VNU_6 VNU61	(.Q1(Q[109])	,.Q2(Q[487])	,.Q3(Q[642])	,.Q4(Q[1014])	,.Q5(Q[1189])	,.Q6(Q[1602])	,.R1(R[109])	,.R2(R[487])	,.R3(R[642])	,.R4(R[1014])	,.R5(R[1189])	,.R6(R[1602])	,.clk(clk)	,.L(L61)	,.P(P[60])	,.reset(reset)	);
VNU_6 VNU62	(.Q1(Q[115])	,.Q2(Q[493])	,.Q3(Q[648])	,.Q4(Q[1020])	,.Q5(Q[1195])	,.Q6(Q[1608])	,.R1(R[115])	,.R2(R[493])	,.R3(R[648])	,.R4(R[1020])	,.R5(R[1195])	,.R6(R[1608])	,.clk(clk)	,.L(L62)	,.P(P[61])	,.reset(reset)	);
VNU_6 VNU63	(.Q1(Q[121])	,.Q2(Q[499])	,.Q3(Q[654])	,.Q4(Q[1026])	,.Q5(Q[1201])	,.Q6(Q[1614])	,.R1(R[121])	,.R2(R[499])	,.R3(R[654])	,.R4(R[1026])	,.R5(R[1201])	,.R6(R[1614])	,.clk(clk)	,.L(L63)	,.P(P[62])	,.reset(reset)	);
VNU_6 VNU64	(.Q1(Q[127])	,.Q2(Q[505])	,.Q3(Q[660])	,.Q4(Q[1032])	,.Q5(Q[1207])	,.Q6(Q[1620])	,.R1(R[127])	,.R2(R[505])	,.R3(R[660])	,.R4(R[1032])	,.R5(R[1207])	,.R6(R[1620])	,.clk(clk)	,.L(L64)	,.P(P[63])	,.reset(reset)	);
VNU_6 VNU65	(.Q1(Q[133])	,.Q2(Q[511])	,.Q3(Q[666])	,.Q4(Q[1038])	,.Q5(Q[1213])	,.Q6(Q[1626])	,.R1(R[133])	,.R2(R[511])	,.R3(R[666])	,.R4(R[1038])	,.R5(R[1213])	,.R6(R[1626])	,.clk(clk)	,.L(L65)	,.P(P[64])	,.reset(reset)	);
VNU_6 VNU66	(.Q1(Q[139])	,.Q2(Q[517])	,.Q3(Q[672])	,.Q4(Q[1044])	,.Q5(Q[1219])	,.Q6(Q[1632])	,.R1(R[139])	,.R2(R[517])	,.R3(R[672])	,.R4(R[1044])	,.R5(R[1219])	,.R6(R[1632])	,.clk(clk)	,.L(L66)	,.P(P[65])	,.reset(reset)	);
VNU_6 VNU67	(.Q1(Q[1])	,.Q2(Q[523])	,.Q3(Q[678])	,.Q4(Q[1050])	,.Q5(Q[1081])	,.Q6(Q[1638])	,.R1(R[1])	,.R2(R[523])	,.R3(R[678])	,.R4(R[1050])	,.R5(R[1081])	,.R6(R[1638])	,.clk(clk)	,.L(L67)	,.P(P[66])	,.reset(reset)	);
VNU_6 VNU68	(.Q1(Q[7])	,.Q2(Q[529])	,.Q3(Q[684])	,.Q4(Q[1056])	,.Q5(Q[1087])	,.Q6(Q[1644])	,.R1(R[7])	,.R2(R[529])	,.R3(R[684])	,.R4(R[1056])	,.R5(R[1087])	,.R6(R[1644])	,.clk(clk)	,.L(L68)	,.P(P[67])	,.reset(reset)	);
VNU_6 VNU69	(.Q1(Q[13])	,.Q2(Q[535])	,.Q3(Q[690])	,.Q4(Q[1062])	,.Q5(Q[1093])	,.Q6(Q[1650])	,.R1(R[13])	,.R2(R[535])	,.R3(R[690])	,.R4(R[1062])	,.R5(R[1093])	,.R6(R[1650])	,.clk(clk)	,.L(L69)	,.P(P[68])	,.reset(reset)	);
VNU_6 VNU70	(.Q1(Q[19])	,.Q2(Q[541])	,.Q3(Q[696])	,.Q4(Q[1068])	,.Q5(Q[1099])	,.Q6(Q[1656])	,.R1(R[19])	,.R2(R[541])	,.R3(R[696])	,.R4(R[1068])	,.R5(R[1099])	,.R6(R[1656])	,.clk(clk)	,.L(L70)	,.P(P[69])	,.reset(reset)	);
VNU_6 VNU71	(.Q1(Q[25])	,.Q2(Q[547])	,.Q3(Q[702])	,.Q4(Q[1074])	,.Q5(Q[1105])	,.Q6(Q[1662])	,.R1(R[25])	,.R2(R[547])	,.R3(R[702])	,.R4(R[1074])	,.R5(R[1105])	,.R6(R[1662])	,.clk(clk)	,.L(L71)	,.P(P[70])	,.reset(reset)	);
VNU_6 VNU72	(.Q1(Q[31])	,.Q2(Q[553])	,.Q3(Q[708])	,.Q4(Q[936])	,.Q5(Q[1111])	,.Q6(Q[1668])	,.R1(R[31])	,.R2(R[553])	,.R3(R[708])	,.R4(R[936])	,.R5(R[1111])	,.R6(R[1668])	,.clk(clk)	,.L(L72)	,.P(P[71])	,.reset(reset)	);
VNU_3 VNU73	(.Q1(Q[438])	,.Q2(Q[1003])	,.Q3(Q[1585])							,.R1(R[438])	,.R2(R[1003])	,.R3(R[1585])							,.clk(clk)	,.L(L73)	,.P(P[72])	,.reset(reset)	);
VNU_3 VNU74	(.Q1(Q[445])	,.Q2(Q[1009])	,.Q3(Q[1591])							,.R1(R[445])	,.R2(R[1009])	,.R3(R[1591])							,.clk(clk)	,.L(L74)	,.P(P[73])	,.reset(reset)	);
VNU_3 VNU75	(.Q1(Q[452])	,.Q2(Q[1015])	,.Q3(Q[1597])							,.R1(R[452])	,.R2(R[1015])	,.R3(R[1597])							,.clk(clk)	,.L(L75)	,.P(P[74])	,.reset(reset)	);
VNU_3 VNU76	(.Q1(Q[459])	,.Q2(Q[1021])	,.Q3(Q[1603])							,.R1(R[459])	,.R2(R[1021])	,.R3(R[1603])							,.clk(clk)	,.L(L76)	,.P(P[75])	,.reset(reset)	);
VNU_3 VNU77	(.Q1(Q[466])	,.Q2(Q[1027])	,.Q3(Q[1609])							,.R1(R[466])	,.R2(R[1027])	,.R3(R[1609])							,.clk(clk)	,.L(L77)	,.P(P[76])	,.reset(reset)	);
VNU_3 VNU78	(.Q1(Q[473])	,.Q2(Q[1033])	,.Q3(Q[1615])							,.R1(R[473])	,.R2(R[1033])	,.R3(R[1615])							,.clk(clk)	,.L(L78)	,.P(P[77])	,.reset(reset)	);
VNU_3 VNU79	(.Q1(Q[312])	,.Q2(Q[1039])	,.Q3(Q[1621])							,.R1(R[312])	,.R2(R[1039])	,.R3(R[1621])							,.clk(clk)	,.L(L79)	,.P(P[78])	,.reset(reset)	);
VNU_3 VNU80	(.Q1(Q[319])	,.Q2(Q[1045])	,.Q3(Q[1627])							,.R1(R[319])	,.R2(R[1045])	,.R3(R[1627])							,.clk(clk)	,.L(L80)	,.P(P[79])	,.reset(reset)	);
VNU_3 VNU81	(.Q1(Q[326])	,.Q2(Q[1051])	,.Q3(Q[1633])							,.R1(R[326])	,.R2(R[1051])	,.R3(R[1633])							,.clk(clk)	,.L(L81)	,.P(P[80])	,.reset(reset)	);
VNU_3 VNU82	(.Q1(Q[333])	,.Q2(Q[1057])	,.Q3(Q[1639])							,.R1(R[333])	,.R2(R[1057])	,.R3(R[1639])							,.clk(clk)	,.L(L82)	,.P(P[81])	,.reset(reset)	);
VNU_3 VNU83	(.Q1(Q[340])	,.Q2(Q[1063])	,.Q3(Q[1645])							,.R1(R[340])	,.R2(R[1063])	,.R3(R[1645])							,.clk(clk)	,.L(L83)	,.P(P[82])	,.reset(reset)	);
VNU_3 VNU84	(.Q1(Q[347])	,.Q2(Q[1069])	,.Q3(Q[1651])							,.R1(R[347])	,.R2(R[1069])	,.R3(R[1651])							,.clk(clk)	,.L(L84)	,.P(P[83])	,.reset(reset)	);
VNU_3 VNU85	(.Q1(Q[354])	,.Q2(Q[1075])	,.Q3(Q[1657])							,.R1(R[354])	,.R2(R[1075])	,.R3(R[1657])							,.clk(clk)	,.L(L85)	,.P(P[84])	,.reset(reset)	);
VNU_3 VNU86	(.Q1(Q[361])	,.Q2(Q[937])	,.Q3(Q[1663])							,.R1(R[361])	,.R2(R[937])	,.R3(R[1663])							,.clk(clk)	,.L(L86)	,.P(P[85])	,.reset(reset)	);
VNU_3 VNU87	(.Q1(Q[368])	,.Q2(Q[943])	,.Q3(Q[1669])							,.R1(R[368])	,.R2(R[943])	,.R3(R[1669])							,.clk(clk)	,.L(L87)	,.P(P[86])	,.reset(reset)	);
VNU_3 VNU88	(.Q1(Q[375])	,.Q2(Q[949])	,.Q3(Q[1675])							,.R1(R[375])	,.R2(R[949])	,.R3(R[1675])							,.clk(clk)	,.L(L88)	,.P(P[87])	,.reset(reset)	);
VNU_3 VNU89	(.Q1(Q[382])	,.Q2(Q[955])	,.Q3(Q[1537])							,.R1(R[382])	,.R2(R[955])	,.R3(R[1537])							,.clk(clk)	,.L(L89)	,.P(P[88])	,.reset(reset)	);
VNU_3 VNU90	(.Q1(Q[389])	,.Q2(Q[961])	,.Q3(Q[1543])							,.R1(R[389])	,.R2(R[961])	,.R3(R[1543])							,.clk(clk)	,.L(L90)	,.P(P[89])	,.reset(reset)	);
VNU_3 VNU91	(.Q1(Q[396])	,.Q2(Q[967])	,.Q3(Q[1549])							,.R1(R[396])	,.R2(R[967])	,.R3(R[1549])							,.clk(clk)	,.L(L91)	,.P(P[90])	,.reset(reset)	);
VNU_3 VNU92	(.Q1(Q[403])	,.Q2(Q[973])	,.Q3(Q[1555])							,.R1(R[403])	,.R2(R[973])	,.R3(R[1555])							,.clk(clk)	,.L(L92)	,.P(P[91])	,.reset(reset)	);
VNU_3 VNU93	(.Q1(Q[410])	,.Q2(Q[979])	,.Q3(Q[1561])							,.R1(R[410])	,.R2(R[979])	,.R3(R[1561])							,.clk(clk)	,.L(L93)	,.P(P[92])	,.reset(reset)	);
VNU_3 VNU94	(.Q1(Q[417])	,.Q2(Q[985])	,.Q3(Q[1567])							,.R1(R[417])	,.R2(R[985])	,.R3(R[1567])							,.clk(clk)	,.L(L94)	,.P(P[93])	,.reset(reset)	);
VNU_3 VNU95	(.Q1(Q[424])	,.Q2(Q[991])	,.Q3(Q[1573])							,.R1(R[424])	,.R2(R[991])	,.R3(R[1573])							,.clk(clk)	,.L(L95)	,.P(P[94])	,.reset(reset)	);
VNU_3 VNU96	(.Q1(Q[431])	,.Q2(Q[997])	,.Q3(Q[1579])							,.R1(R[431])	,.R2(R[997])	,.R3(R[1579])							,.clk(clk)	,.L(L96)	,.P(P[95])	,.reset(reset)	);
VNU_3 VNU97	(.Q1(Q[446])	,.Q2(Q[859])	,.Q3(Q[1253])							,.R1(R[446])	,.R2(R[859])	,.R3(R[1253])							,.clk(clk)	,.L(L97)	,.P(P[96])	,.reset(reset)	);
VNU_3 VNU98	(.Q1(Q[453])	,.Q2(Q[866])	,.Q3(Q[1260])							,.R1(R[453])	,.R2(R[866])	,.R3(R[1260])							,.clk(clk)	,.L(L98)	,.P(P[97])	,.reset(reset)	);
VNU_3 VNU99	(.Q1(Q[460])	,.Q2(Q[873])	,.Q3(Q[1267])							,.R1(R[460])	,.R2(R[873])	,.R3(R[1267])							,.clk(clk)	,.L(L99)	,.P(P[98])	,.reset(reset)	);
VNU_3 VNU100	(.Q1(Q[467])	,.Q2(Q[880])	,.Q3(Q[1274])							,.R1(R[467])	,.R2(R[880])	,.R3(R[1274])							,.clk(clk)	,.L(L100)	,.P(P[99])	,.reset(reset)	);
VNU_3 VNU101	(.Q1(Q[474])	,.Q2(Q[887])	,.Q3(Q[1281])							,.R1(R[474])	,.R2(R[887])	,.R3(R[1281])							,.clk(clk)	,.L(L101)	,.P(P[100])	,.reset(reset)	);
VNU_3 VNU102	(.Q1(Q[313])	,.Q2(Q[894])	,.Q3(Q[1288])							,.R1(R[313])	,.R2(R[894])	,.R3(R[1288])							,.clk(clk)	,.L(L102)	,.P(P[101])	,.reset(reset)	);
VNU_3 VNU103	(.Q1(Q[320])	,.Q2(Q[901])	,.Q3(Q[1295])							,.R1(R[320])	,.R2(R[901])	,.R3(R[1295])							,.clk(clk)	,.L(L103)	,.P(P[102])	,.reset(reset)	);
VNU_3 VNU104	(.Q1(Q[327])	,.Q2(Q[908])	,.Q3(Q[1302])							,.R1(R[327])	,.R2(R[908])	,.R3(R[1302])							,.clk(clk)	,.L(L104)	,.P(P[103])	,.reset(reset)	);
VNU_3 VNU105	(.Q1(Q[334])	,.Q2(Q[915])	,.Q3(Q[1309])							,.R1(R[334])	,.R2(R[915])	,.R3(R[1309])							,.clk(clk)	,.L(L105)	,.P(P[104])	,.reset(reset)	);
VNU_3 VNU106	(.Q1(Q[341])	,.Q2(Q[922])	,.Q3(Q[1316])							,.R1(R[341])	,.R2(R[922])	,.R3(R[1316])							,.clk(clk)	,.L(L106)	,.P(P[105])	,.reset(reset)	);
VNU_3 VNU107	(.Q1(Q[348])	,.Q2(Q[929])	,.Q3(Q[1323])							,.R1(R[348])	,.R2(R[929])	,.R3(R[1323])							,.clk(clk)	,.L(L107)	,.P(P[106])	,.reset(reset)	);
VNU_3 VNU108	(.Q1(Q[355])	,.Q2(Q[768])	,.Q3(Q[1330])							,.R1(R[355])	,.R2(R[768])	,.R3(R[1330])							,.clk(clk)	,.L(L108)	,.P(P[107])	,.reset(reset)	);
VNU_3 VNU109	(.Q1(Q[362])	,.Q2(Q[775])	,.Q3(Q[1337])							,.R1(R[362])	,.R2(R[775])	,.R3(R[1337])							,.clk(clk)	,.L(L109)	,.P(P[108])	,.reset(reset)	);
VNU_3 VNU110	(.Q1(Q[369])	,.Q2(Q[782])	,.Q3(Q[1344])							,.R1(R[369])	,.R2(R[782])	,.R3(R[1344])							,.clk(clk)	,.L(L110)	,.P(P[109])	,.reset(reset)	);
VNU_3 VNU111	(.Q1(Q[376])	,.Q2(Q[789])	,.Q3(Q[1351])							,.R1(R[376])	,.R2(R[789])	,.R3(R[1351])							,.clk(clk)	,.L(L111)	,.P(P[110])	,.reset(reset)	);
VNU_3 VNU112	(.Q1(Q[383])	,.Q2(Q[796])	,.Q3(Q[1358])							,.R1(R[383])	,.R2(R[796])	,.R3(R[1358])							,.clk(clk)	,.L(L112)	,.P(P[111])	,.reset(reset)	);
VNU_3 VNU113	(.Q1(Q[390])	,.Q2(Q[803])	,.Q3(Q[1365])							,.R1(R[390])	,.R2(R[803])	,.R3(R[1365])							,.clk(clk)	,.L(L113)	,.P(P[112])	,.reset(reset)	);
VNU_3 VNU114	(.Q1(Q[397])	,.Q2(Q[810])	,.Q3(Q[1372])							,.R1(R[397])	,.R2(R[810])	,.R3(R[1372])							,.clk(clk)	,.L(L114)	,.P(P[113])	,.reset(reset)	);
VNU_3 VNU115	(.Q1(Q[404])	,.Q2(Q[817])	,.Q3(Q[1379])							,.R1(R[404])	,.R2(R[817])	,.R3(R[1379])							,.clk(clk)	,.L(L115)	,.P(P[114])	,.reset(reset)	);
VNU_3 VNU116	(.Q1(Q[411])	,.Q2(Q[824])	,.Q3(Q[1386])							,.R1(R[411])	,.R2(R[824])	,.R3(R[1386])							,.clk(clk)	,.L(L116)	,.P(P[115])	,.reset(reset)	);
VNU_3 VNU117	(.Q1(Q[418])	,.Q2(Q[831])	,.Q3(Q[1225])							,.R1(R[418])	,.R2(R[831])	,.R3(R[1225])							,.clk(clk)	,.L(L117)	,.P(P[116])	,.reset(reset)	);
VNU_3 VNU118	(.Q1(Q[425])	,.Q2(Q[838])	,.Q3(Q[1232])							,.R1(R[425])	,.R2(R[838])	,.R3(R[1232])							,.clk(clk)	,.L(L118)	,.P(P[117])	,.reset(reset)	);
VNU_3 VNU119	(.Q1(Q[432])	,.Q2(Q[845])	,.Q3(Q[1239])							,.R1(R[432])	,.R2(R[845])	,.R3(R[1239])							,.clk(clk)	,.L(L119)	,.P(P[118])	,.reset(reset)	);
VNU_3 VNU120	(.Q1(Q[439])	,.Q2(Q[852])	,.Q3(Q[1246])							,.R1(R[439])	,.R2(R[852])	,.R3(R[1246])							,.clk(clk)	,.L(L120)	,.P(P[119])	,.reset(reset)	);
VNU_6 VNU121	(.Q1(Q[278])	,.Q2(Q[342])	,.Q3(Q[867])	,.Q4(Q[1352])	,.Q5(Q[1398])	,.Q6(Q[1729])	,.R1(R[278])	,.R2(R[342])	,.R3(R[867])	,.R4(R[1352])	,.R5(R[1398])	,.R6(R[1729])	,.clk(clk)	,.L(L121)	,.P(P[120])	,.reset(reset)	);
VNU_6 VNU122	(.Q1(Q[285])	,.Q2(Q[349])	,.Q3(Q[874])	,.Q4(Q[1359])	,.Q5(Q[1404])	,.Q6(Q[1735])	,.R1(R[285])	,.R2(R[349])	,.R3(R[874])	,.R4(R[1359])	,.R5(R[1404])	,.R6(R[1735])	,.clk(clk)	,.L(L122)	,.P(P[121])	,.reset(reset)	);
VNU_6 VNU123	(.Q1(Q[292])	,.Q2(Q[356])	,.Q3(Q[881])	,.Q4(Q[1366])	,.Q5(Q[1410])	,.Q6(Q[1741])	,.R1(R[292])	,.R2(R[356])	,.R3(R[881])	,.R4(R[1366])	,.R5(R[1410])	,.R6(R[1741])	,.clk(clk)	,.L(L123)	,.P(P[122])	,.reset(reset)	);
VNU_6 VNU124	(.Q1(Q[299])	,.Q2(Q[363])	,.Q3(Q[888])	,.Q4(Q[1373])	,.Q5(Q[1416])	,.Q6(Q[1747])	,.R1(R[299])	,.R2(R[363])	,.R3(R[888])	,.R4(R[1373])	,.R5(R[1416])	,.R6(R[1747])	,.clk(clk)	,.L(L124)	,.P(P[123])	,.reset(reset)	);
VNU_6 VNU125	(.Q1(Q[306])	,.Q2(Q[370])	,.Q3(Q[895])	,.Q4(Q[1380])	,.Q5(Q[1422])	,.Q6(Q[1753])	,.R1(R[306])	,.R2(R[370])	,.R3(R[895])	,.R4(R[1380])	,.R5(R[1422])	,.R6(R[1753])	,.clk(clk)	,.L(L125)	,.P(P[124])	,.reset(reset)	);
VNU_6 VNU126	(.Q1(Q[145])	,.Q2(Q[377])	,.Q3(Q[902])	,.Q4(Q[1387])	,.Q5(Q[1428])	,.Q6(Q[1759])	,.R1(R[145])	,.R2(R[377])	,.R3(R[902])	,.R4(R[1387])	,.R5(R[1428])	,.R6(R[1759])	,.clk(clk)	,.L(L126)	,.P(P[125])	,.reset(reset)	);
VNU_6 VNU127	(.Q1(Q[152])	,.Q2(Q[384])	,.Q3(Q[909])	,.Q4(Q[1226])	,.Q5(Q[1434])	,.Q6(Q[1765])	,.R1(R[152])	,.R2(R[384])	,.R3(R[909])	,.R4(R[1226])	,.R5(R[1434])	,.R6(R[1765])	,.clk(clk)	,.L(L127)	,.P(P[126])	,.reset(reset)	);
VNU_6 VNU128	(.Q1(Q[159])	,.Q2(Q[391])	,.Q3(Q[916])	,.Q4(Q[1233])	,.Q5(Q[1440])	,.Q6(Q[1771])	,.R1(R[159])	,.R2(R[391])	,.R3(R[916])	,.R4(R[1233])	,.R5(R[1440])	,.R6(R[1771])	,.clk(clk)	,.L(L128)	,.P(P[127])	,.reset(reset)	);
VNU_6 VNU129	(.Q1(Q[166])	,.Q2(Q[398])	,.Q3(Q[923])	,.Q4(Q[1240])	,.Q5(Q[1446])	,.Q6(Q[1777])	,.R1(R[166])	,.R2(R[398])	,.R3(R[923])	,.R4(R[1240])	,.R5(R[1446])	,.R6(R[1777])	,.clk(clk)	,.L(L129)	,.P(P[128])	,.reset(reset)	);
VNU_6 VNU130	(.Q1(Q[173])	,.Q2(Q[405])	,.Q3(Q[930])	,.Q4(Q[1247])	,.Q5(Q[1452])	,.Q6(Q[1783])	,.R1(R[173])	,.R2(R[405])	,.R3(R[930])	,.R4(R[1247])	,.R5(R[1452])	,.R6(R[1783])	,.clk(clk)	,.L(L130)	,.P(P[129])	,.reset(reset)	);
VNU_6 VNU131	(.Q1(Q[180])	,.Q2(Q[412])	,.Q3(Q[769])	,.Q4(Q[1254])	,.Q5(Q[1458])	,.Q6(Q[1789])	,.R1(R[180])	,.R2(R[412])	,.R3(R[769])	,.R4(R[1254])	,.R5(R[1458])	,.R6(R[1789])	,.clk(clk)	,.L(L131)	,.P(P[130])	,.reset(reset)	);
VNU_6 VNU132	(.Q1(Q[187])	,.Q2(Q[419])	,.Q3(Q[776])	,.Q4(Q[1261])	,.Q5(Q[1464])	,.Q6(Q[1795])	,.R1(R[187])	,.R2(R[419])	,.R3(R[776])	,.R4(R[1261])	,.R5(R[1464])	,.R6(R[1795])	,.clk(clk)	,.L(L132)	,.P(P[131])	,.reset(reset)	);
VNU_6 VNU133	(.Q1(Q[194])	,.Q2(Q[426])	,.Q3(Q[783])	,.Q4(Q[1268])	,.Q5(Q[1470])	,.Q6(Q[1801])	,.R1(R[194])	,.R2(R[426])	,.R3(R[783])	,.R4(R[1268])	,.R5(R[1470])	,.R6(R[1801])	,.clk(clk)	,.L(L133)	,.P(P[132])	,.reset(reset)	);
VNU_6 VNU134	(.Q1(Q[201])	,.Q2(Q[433])	,.Q3(Q[790])	,.Q4(Q[1275])	,.Q5(Q[1476])	,.Q6(Q[1807])	,.R1(R[201])	,.R2(R[433])	,.R3(R[790])	,.R4(R[1275])	,.R5(R[1476])	,.R6(R[1807])	,.clk(clk)	,.L(L134)	,.P(P[133])	,.reset(reset)	);
VNU_6 VNU135	(.Q1(Q[208])	,.Q2(Q[440])	,.Q3(Q[797])	,.Q4(Q[1282])	,.Q5(Q[1482])	,.Q6(Q[1813])	,.R1(R[208])	,.R2(R[440])	,.R3(R[797])	,.R4(R[1282])	,.R5(R[1482])	,.R6(R[1813])	,.clk(clk)	,.L(L135)	,.P(P[134])	,.reset(reset)	);
VNU_6 VNU136	(.Q1(Q[215])	,.Q2(Q[447])	,.Q3(Q[804])	,.Q4(Q[1289])	,.Q5(Q[1488])	,.Q6(Q[1819])	,.R1(R[215])	,.R2(R[447])	,.R3(R[804])	,.R4(R[1289])	,.R5(R[1488])	,.R6(R[1819])	,.clk(clk)	,.L(L136)	,.P(P[135])	,.reset(reset)	);
VNU_6 VNU137	(.Q1(Q[222])	,.Q2(Q[454])	,.Q3(Q[811])	,.Q4(Q[1296])	,.Q5(Q[1494])	,.Q6(Q[1681])	,.R1(R[222])	,.R2(R[454])	,.R3(R[811])	,.R4(R[1296])	,.R5(R[1494])	,.R6(R[1681])	,.clk(clk)	,.L(L137)	,.P(P[136])	,.reset(reset)	);
VNU_6 VNU138	(.Q1(Q[229])	,.Q2(Q[461])	,.Q3(Q[818])	,.Q4(Q[1303])	,.Q5(Q[1500])	,.Q6(Q[1687])	,.R1(R[229])	,.R2(R[461])	,.R3(R[818])	,.R4(R[1303])	,.R5(R[1500])	,.R6(R[1687])	,.clk(clk)	,.L(L138)	,.P(P[137])	,.reset(reset)	);
VNU_6 VNU139	(.Q1(Q[236])	,.Q2(Q[468])	,.Q3(Q[825])	,.Q4(Q[1310])	,.Q5(Q[1506])	,.Q6(Q[1693])	,.R1(R[236])	,.R2(R[468])	,.R3(R[825])	,.R4(R[1310])	,.R5(R[1506])	,.R6(R[1693])	,.clk(clk)	,.L(L139)	,.P(P[138])	,.reset(reset)	);
VNU_6 VNU140	(.Q1(Q[243])	,.Q2(Q[475])	,.Q3(Q[832])	,.Q4(Q[1317])	,.Q5(Q[1512])	,.Q6(Q[1699])	,.R1(R[243])	,.R2(R[475])	,.R3(R[832])	,.R4(R[1317])	,.R5(R[1512])	,.R6(R[1699])	,.clk(clk)	,.L(L140)	,.P(P[139])	,.reset(reset)	);
VNU_6 VNU141	(.Q1(Q[250])	,.Q2(Q[314])	,.Q3(Q[839])	,.Q4(Q[1324])	,.Q5(Q[1518])	,.Q6(Q[1705])	,.R1(R[250])	,.R2(R[314])	,.R3(R[839])	,.R4(R[1324])	,.R5(R[1518])	,.R6(R[1705])	,.clk(clk)	,.L(L141)	,.P(P[140])	,.reset(reset)	);
VNU_6 VNU142	(.Q1(Q[257])	,.Q2(Q[321])	,.Q3(Q[846])	,.Q4(Q[1331])	,.Q5(Q[1524])	,.Q6(Q[1711])	,.R1(R[257])	,.R2(R[321])	,.R3(R[846])	,.R4(R[1331])	,.R5(R[1524])	,.R6(R[1711])	,.clk(clk)	,.L(L142)	,.P(P[141])	,.reset(reset)	);
VNU_6 VNU143	(.Q1(Q[264])	,.Q2(Q[328])	,.Q3(Q[853])	,.Q4(Q[1338])	,.Q5(Q[1530])	,.Q6(Q[1717])	,.R1(R[264])	,.R2(R[328])	,.R3(R[853])	,.R4(R[1338])	,.R5(R[1530])	,.R6(R[1717])	,.clk(clk)	,.L(L143)	,.P(P[142])	,.reset(reset)	);
VNU_6 VNU144	(.Q1(Q[271])	,.Q2(Q[335])	,.Q3(Q[860])	,.Q4(Q[1345])	,.Q5(Q[1392])	,.Q6(Q[1723])	,.R1(R[271])	,.R2(R[335])	,.R3(R[860])	,.R4(R[1345])	,.R5(R[1392])	,.R6(R[1723])	,.clk(clk)	,.L(L144)	,.P(P[143])	,.reset(reset)	);
VNU_3 VNU145	(.Q1(Q[181])	,.Q2(Q[643])	,.Q3(Q[1082])							,.R1(R[181])	,.R2(R[643])	,.R3(R[1082])							,.clk(clk)	,.L(L145)	,.P(P[144])	,.reset(reset)	);
VNU_3 VNU146	(.Q1(Q[188])	,.Q2(Q[649])	,.Q3(Q[1088])							,.R1(R[188])	,.R2(R[649])	,.R3(R[1088])							,.clk(clk)	,.L(L146)	,.P(P[145])	,.reset(reset)	);
VNU_3 VNU147	(.Q1(Q[195])	,.Q2(Q[655])	,.Q3(Q[1094])							,.R1(R[195])	,.R2(R[655])	,.R3(R[1094])							,.clk(clk)	,.L(L147)	,.P(P[146])	,.reset(reset)	);
VNU_3 VNU148	(.Q1(Q[202])	,.Q2(Q[661])	,.Q3(Q[1100])							,.R1(R[202])	,.R2(R[661])	,.R3(R[1100])							,.clk(clk)	,.L(L148)	,.P(P[147])	,.reset(reset)	);
VNU_3 VNU149	(.Q1(Q[209])	,.Q2(Q[667])	,.Q3(Q[1106])							,.R1(R[209])	,.R2(R[667])	,.R3(R[1106])							,.clk(clk)	,.L(L149)	,.P(P[148])	,.reset(reset)	);
VNU_3 VNU150	(.Q1(Q[216])	,.Q2(Q[673])	,.Q3(Q[1112])							,.R1(R[216])	,.R2(R[673])	,.R3(R[1112])							,.clk(clk)	,.L(L150)	,.P(P[149])	,.reset(reset)	);
VNU_3 VNU151	(.Q1(Q[223])	,.Q2(Q[679])	,.Q3(Q[1118])							,.R1(R[223])	,.R2(R[679])	,.R3(R[1118])							,.clk(clk)	,.L(L151)	,.P(P[150])	,.reset(reset)	);
VNU_3 VNU152	(.Q1(Q[230])	,.Q2(Q[685])	,.Q3(Q[1124])							,.R1(R[230])	,.R2(R[685])	,.R3(R[1124])							,.clk(clk)	,.L(L152)	,.P(P[151])	,.reset(reset)	);
VNU_3 VNU153	(.Q1(Q[237])	,.Q2(Q[691])	,.Q3(Q[1130])							,.R1(R[237])	,.R2(R[691])	,.R3(R[1130])							,.clk(clk)	,.L(L153)	,.P(P[152])	,.reset(reset)	);
VNU_3 VNU154	(.Q1(Q[244])	,.Q2(Q[697])	,.Q3(Q[1136])							,.R1(R[244])	,.R2(R[697])	,.R3(R[1136])							,.clk(clk)	,.L(L154)	,.P(P[153])	,.reset(reset)	);
VNU_3 VNU155	(.Q1(Q[251])	,.Q2(Q[703])	,.Q3(Q[1142])							,.R1(R[251])	,.R2(R[703])	,.R3(R[1142])							,.clk(clk)	,.L(L155)	,.P(P[154])	,.reset(reset)	);
VNU_3 VNU156	(.Q1(Q[258])	,.Q2(Q[709])	,.Q3(Q[1148])							,.R1(R[258])	,.R2(R[709])	,.R3(R[1148])							,.clk(clk)	,.L(L156)	,.P(P[155])	,.reset(reset)	);
VNU_3 VNU157	(.Q1(Q[265])	,.Q2(Q[715])	,.Q3(Q[1154])							,.R1(R[265])	,.R2(R[715])	,.R3(R[1154])							,.clk(clk)	,.L(L157)	,.P(P[156])	,.reset(reset)	);
VNU_3 VNU158	(.Q1(Q[272])	,.Q2(Q[721])	,.Q3(Q[1160])							,.R1(R[272])	,.R2(R[721])	,.R3(R[1160])							,.clk(clk)	,.L(L158)	,.P(P[157])	,.reset(reset)	);
VNU_3 VNU159	(.Q1(Q[279])	,.Q2(Q[727])	,.Q3(Q[1166])							,.R1(R[279])	,.R2(R[727])	,.R3(R[1166])							,.clk(clk)	,.L(L159)	,.P(P[158])	,.reset(reset)	);
VNU_3 VNU160	(.Q1(Q[286])	,.Q2(Q[733])	,.Q3(Q[1172])							,.R1(R[286])	,.R2(R[733])	,.R3(R[1172])							,.clk(clk)	,.L(L160)	,.P(P[159])	,.reset(reset)	);
VNU_3 VNU161	(.Q1(Q[293])	,.Q2(Q[739])	,.Q3(Q[1178])							,.R1(R[293])	,.R2(R[739])	,.R3(R[1178])							,.clk(clk)	,.L(L161)	,.P(P[160])	,.reset(reset)	);
VNU_3 VNU162	(.Q1(Q[300])	,.Q2(Q[745])	,.Q3(Q[1184])							,.R1(R[300])	,.R2(R[745])	,.R3(R[1184])							,.clk(clk)	,.L(L162)	,.P(P[161])	,.reset(reset)	);
VNU_3 VNU163	(.Q1(Q[307])	,.Q2(Q[751])	,.Q3(Q[1190])							,.R1(R[307])	,.R2(R[751])	,.R3(R[1190])							,.clk(clk)	,.L(L163)	,.P(P[162])	,.reset(reset)	);
VNU_3 VNU164	(.Q1(Q[146])	,.Q2(Q[757])	,.Q3(Q[1196])							,.R1(R[146])	,.R2(R[757])	,.R3(R[1196])							,.clk(clk)	,.L(L164)	,.P(P[163])	,.reset(reset)	);
VNU_3 VNU165	(.Q1(Q[153])	,.Q2(Q[763])	,.Q3(Q[1202])							,.R1(R[153])	,.R2(R[763])	,.R3(R[1202])							,.clk(clk)	,.L(L165)	,.P(P[164])	,.reset(reset)	);
VNU_3 VNU166	(.Q1(Q[160])	,.Q2(Q[625])	,.Q3(Q[1208])							,.R1(R[160])	,.R2(R[625])	,.R3(R[1208])							,.clk(clk)	,.L(L166)	,.P(P[165])	,.reset(reset)	);
VNU_3 VNU167	(.Q1(Q[167])	,.Q2(Q[631])	,.Q3(Q[1214])							,.R1(R[167])	,.R2(R[631])	,.R3(R[1214])							,.clk(clk)	,.L(L167)	,.P(P[166])	,.reset(reset)	);
VNU_3 VNU168	(.Q1(Q[174])	,.Q2(Q[637])	,.Q3(Q[1220])							,.R1(R[174])	,.R2(R[637])	,.R3(R[1220])							,.clk(clk)	,.L(L168)	,.P(P[167])	,.reset(reset)	);
VNU_6 VNU169	(.Q1(Q[301])	,.Q2(Q[427])	,.Q3(Q[798])	,.Q4(Q[1325])	,.Q5(Q[1453])	,.Q6(Q[1766])	,.R1(R[301])	,.R2(R[427])	,.R3(R[798])	,.R4(R[1325])	,.R5(R[1453])	,.R6(R[1766])	,.clk(clk)	,.L(L169)	,.P(P[168])	,.reset(reset)	);
VNU_6 VNU170	(.Q1(Q[308])	,.Q2(Q[434])	,.Q3(Q[805])	,.Q4(Q[1332])	,.Q5(Q[1459])	,.Q6(Q[1772])	,.R1(R[308])	,.R2(R[434])	,.R3(R[805])	,.R4(R[1332])	,.R5(R[1459])	,.R6(R[1772])	,.clk(clk)	,.L(L170)	,.P(P[169])	,.reset(reset)	);
VNU_6 VNU171	(.Q1(Q[147])	,.Q2(Q[441])	,.Q3(Q[812])	,.Q4(Q[1339])	,.Q5(Q[1465])	,.Q6(Q[1778])	,.R1(R[147])	,.R2(R[441])	,.R3(R[812])	,.R4(R[1339])	,.R5(R[1465])	,.R6(R[1778])	,.clk(clk)	,.L(L171)	,.P(P[170])	,.reset(reset)	);
VNU_6 VNU172	(.Q1(Q[154])	,.Q2(Q[448])	,.Q3(Q[819])	,.Q4(Q[1346])	,.Q5(Q[1471])	,.Q6(Q[1784])	,.R1(R[154])	,.R2(R[448])	,.R3(R[819])	,.R4(R[1346])	,.R5(R[1471])	,.R6(R[1784])	,.clk(clk)	,.L(L172)	,.P(P[171])	,.reset(reset)	);
VNU_6 VNU173	(.Q1(Q[161])	,.Q2(Q[455])	,.Q3(Q[826])	,.Q4(Q[1353])	,.Q5(Q[1477])	,.Q6(Q[1790])	,.R1(R[161])	,.R2(R[455])	,.R3(R[826])	,.R4(R[1353])	,.R5(R[1477])	,.R6(R[1790])	,.clk(clk)	,.L(L173)	,.P(P[172])	,.reset(reset)	);
VNU_6 VNU174	(.Q1(Q[168])	,.Q2(Q[462])	,.Q3(Q[833])	,.Q4(Q[1360])	,.Q5(Q[1483])	,.Q6(Q[1796])	,.R1(R[168])	,.R2(R[462])	,.R3(R[833])	,.R4(R[1360])	,.R5(R[1483])	,.R6(R[1796])	,.clk(clk)	,.L(L174)	,.P(P[173])	,.reset(reset)	);
VNU_6 VNU175	(.Q1(Q[175])	,.Q2(Q[469])	,.Q3(Q[840])	,.Q4(Q[1367])	,.Q5(Q[1489])	,.Q6(Q[1802])	,.R1(R[175])	,.R2(R[469])	,.R3(R[840])	,.R4(R[1367])	,.R5(R[1489])	,.R6(R[1802])	,.clk(clk)	,.L(L175)	,.P(P[174])	,.reset(reset)	);
VNU_6 VNU176	(.Q1(Q[182])	,.Q2(Q[476])	,.Q3(Q[847])	,.Q4(Q[1374])	,.Q5(Q[1495])	,.Q6(Q[1808])	,.R1(R[182])	,.R2(R[476])	,.R3(R[847])	,.R4(R[1374])	,.R5(R[1495])	,.R6(R[1808])	,.clk(clk)	,.L(L176)	,.P(P[175])	,.reset(reset)	);
VNU_6 VNU177	(.Q1(Q[189])	,.Q2(Q[315])	,.Q3(Q[854])	,.Q4(Q[1381])	,.Q5(Q[1501])	,.Q6(Q[1814])	,.R1(R[189])	,.R2(R[315])	,.R3(R[854])	,.R4(R[1381])	,.R5(R[1501])	,.R6(R[1814])	,.clk(clk)	,.L(L177)	,.P(P[176])	,.reset(reset)	);
VNU_6 VNU178	(.Q1(Q[196])	,.Q2(Q[322])	,.Q3(Q[861])	,.Q4(Q[1388])	,.Q5(Q[1507])	,.Q6(Q[1820])	,.R1(R[196])	,.R2(R[322])	,.R3(R[861])	,.R4(R[1388])	,.R5(R[1507])	,.R6(R[1820])	,.clk(clk)	,.L(L178)	,.P(P[177])	,.reset(reset)	);
VNU_6 VNU179	(.Q1(Q[203])	,.Q2(Q[329])	,.Q3(Q[868])	,.Q4(Q[1227])	,.Q5(Q[1513])	,.Q6(Q[1682])	,.R1(R[203])	,.R2(R[329])	,.R3(R[868])	,.R4(R[1227])	,.R5(R[1513])	,.R6(R[1682])	,.clk(clk)	,.L(L179)	,.P(P[178])	,.reset(reset)	);
VNU_6 VNU180	(.Q1(Q[210])	,.Q2(Q[336])	,.Q3(Q[875])	,.Q4(Q[1234])	,.Q5(Q[1519])	,.Q6(Q[1688])	,.R1(R[210])	,.R2(R[336])	,.R3(R[875])	,.R4(R[1234])	,.R5(R[1519])	,.R6(R[1688])	,.clk(clk)	,.L(L180)	,.P(P[179])	,.reset(reset)	);
VNU_6 VNU181	(.Q1(Q[217])	,.Q2(Q[343])	,.Q3(Q[882])	,.Q4(Q[1241])	,.Q5(Q[1525])	,.Q6(Q[1694])	,.R1(R[217])	,.R2(R[343])	,.R3(R[882])	,.R4(R[1241])	,.R5(R[1525])	,.R6(R[1694])	,.clk(clk)	,.L(L181)	,.P(P[180])	,.reset(reset)	);
VNU_6 VNU182	(.Q1(Q[224])	,.Q2(Q[350])	,.Q3(Q[889])	,.Q4(Q[1248])	,.Q5(Q[1531])	,.Q6(Q[1700])	,.R1(R[224])	,.R2(R[350])	,.R3(R[889])	,.R4(R[1248])	,.R5(R[1531])	,.R6(R[1700])	,.clk(clk)	,.L(L182)	,.P(P[181])	,.reset(reset)	);
VNU_6 VNU183	(.Q1(Q[231])	,.Q2(Q[357])	,.Q3(Q[896])	,.Q4(Q[1255])	,.Q5(Q[1393])	,.Q6(Q[1706])	,.R1(R[231])	,.R2(R[357])	,.R3(R[896])	,.R4(R[1255])	,.R5(R[1393])	,.R6(R[1706])	,.clk(clk)	,.L(L183)	,.P(P[182])	,.reset(reset)	);
VNU_6 VNU184	(.Q1(Q[238])	,.Q2(Q[364])	,.Q3(Q[903])	,.Q4(Q[1262])	,.Q5(Q[1399])	,.Q6(Q[1712])	,.R1(R[238])	,.R2(R[364])	,.R3(R[903])	,.R4(R[1262])	,.R5(R[1399])	,.R6(R[1712])	,.clk(clk)	,.L(L184)	,.P(P[183])	,.reset(reset)	);
VNU_6 VNU185	(.Q1(Q[245])	,.Q2(Q[371])	,.Q3(Q[910])	,.Q4(Q[1269])	,.Q5(Q[1405])	,.Q6(Q[1718])	,.R1(R[245])	,.R2(R[371])	,.R3(R[910])	,.R4(R[1269])	,.R5(R[1405])	,.R6(R[1718])	,.clk(clk)	,.L(L185)	,.P(P[184])	,.reset(reset)	);
VNU_6 VNU186	(.Q1(Q[252])	,.Q2(Q[378])	,.Q3(Q[917])	,.Q4(Q[1276])	,.Q5(Q[1411])	,.Q6(Q[1724])	,.R1(R[252])	,.R2(R[378])	,.R3(R[917])	,.R4(R[1276])	,.R5(R[1411])	,.R6(R[1724])	,.clk(clk)	,.L(L186)	,.P(P[185])	,.reset(reset)	);
VNU_6 VNU187	(.Q1(Q[259])	,.Q2(Q[385])	,.Q3(Q[924])	,.Q4(Q[1283])	,.Q5(Q[1417])	,.Q6(Q[1730])	,.R1(R[259])	,.R2(R[385])	,.R3(R[924])	,.R4(R[1283])	,.R5(R[1417])	,.R6(R[1730])	,.clk(clk)	,.L(L187)	,.P(P[186])	,.reset(reset)	);
VNU_6 VNU188	(.Q1(Q[266])	,.Q2(Q[392])	,.Q3(Q[931])	,.Q4(Q[1290])	,.Q5(Q[1423])	,.Q6(Q[1736])	,.R1(R[266])	,.R2(R[392])	,.R3(R[931])	,.R4(R[1290])	,.R5(R[1423])	,.R6(R[1736])	,.clk(clk)	,.L(L188)	,.P(P[187])	,.reset(reset)	);
VNU_6 VNU189	(.Q1(Q[273])	,.Q2(Q[399])	,.Q3(Q[770])	,.Q4(Q[1297])	,.Q5(Q[1429])	,.Q6(Q[1742])	,.R1(R[273])	,.R2(R[399])	,.R3(R[770])	,.R4(R[1297])	,.R5(R[1429])	,.R6(R[1742])	,.clk(clk)	,.L(L189)	,.P(P[188])	,.reset(reset)	);
VNU_6 VNU190	(.Q1(Q[280])	,.Q2(Q[406])	,.Q3(Q[777])	,.Q4(Q[1304])	,.Q5(Q[1435])	,.Q6(Q[1748])	,.R1(R[280])	,.R2(R[406])	,.R3(R[777])	,.R4(R[1304])	,.R5(R[1435])	,.R6(R[1748])	,.clk(clk)	,.L(L190)	,.P(P[189])	,.reset(reset)	);
VNU_6 VNU191	(.Q1(Q[287])	,.Q2(Q[413])	,.Q3(Q[784])	,.Q4(Q[1311])	,.Q5(Q[1441])	,.Q6(Q[1754])	,.R1(R[287])	,.R2(R[413])	,.R3(R[784])	,.R4(R[1311])	,.R5(R[1441])	,.R6(R[1754])	,.clk(clk)	,.L(L191)	,.P(P[190])	,.reset(reset)	);
VNU_6 VNU192	(.Q1(Q[294])	,.Q2(Q[420])	,.Q3(Q[791])	,.Q4(Q[1318])	,.Q5(Q[1447])	,.Q6(Q[1760])	,.R1(R[294])	,.R2(R[420])	,.R3(R[791])	,.R4(R[1318])	,.R5(R[1447])	,.R6(R[1760])	,.clk(clk)	,.L(L192)	,.P(P[191])	,.reset(reset)	);
VNU_3 VNU193	(.Q1(Q[68])	,.Q2(Q[530])	,.Q3(Q[1628])							,.R1(R[68])	,.R2(R[530])	,.R3(R[1628])							,.clk(clk)	,.L(L193)	,.P(P[192])	,.reset(reset)	);
VNU_3 VNU194	(.Q1(Q[74])	,.Q2(Q[536])	,.Q3(Q[1634])							,.R1(R[74])	,.R2(R[536])	,.R3(R[1634])							,.clk(clk)	,.L(L194)	,.P(P[193])	,.reset(reset)	);
VNU_3 VNU195	(.Q1(Q[80])	,.Q2(Q[542])	,.Q3(Q[1640])							,.R1(R[80])	,.R2(R[542])	,.R3(R[1640])							,.clk(clk)	,.L(L195)	,.P(P[194])	,.reset(reset)	);
VNU_3 VNU196	(.Q1(Q[86])	,.Q2(Q[548])	,.Q3(Q[1646])							,.R1(R[86])	,.R2(R[548])	,.R3(R[1646])							,.clk(clk)	,.L(L196)	,.P(P[195])	,.reset(reset)	);
VNU_3 VNU197	(.Q1(Q[92])	,.Q2(Q[554])	,.Q3(Q[1652])							,.R1(R[92])	,.R2(R[554])	,.R3(R[1652])							,.clk(clk)	,.L(L197)	,.P(P[196])	,.reset(reset)	);
VNU_3 VNU198	(.Q1(Q[98])	,.Q2(Q[560])	,.Q3(Q[1658])							,.R1(R[98])	,.R2(R[560])	,.R3(R[1658])							,.clk(clk)	,.L(L198)	,.P(P[197])	,.reset(reset)	);
VNU_3 VNU199	(.Q1(Q[104])	,.Q2(Q[566])	,.Q3(Q[1664])							,.R1(R[104])	,.R2(R[566])	,.R3(R[1664])							,.clk(clk)	,.L(L199)	,.P(P[198])	,.reset(reset)	);
VNU_3 VNU200	(.Q1(Q[110])	,.Q2(Q[572])	,.Q3(Q[1670])							,.R1(R[110])	,.R2(R[572])	,.R3(R[1670])							,.clk(clk)	,.L(L200)	,.P(P[199])	,.reset(reset)	);
VNU_3 VNU201	(.Q1(Q[116])	,.Q2(Q[578])	,.Q3(Q[1676])							,.R1(R[116])	,.R2(R[578])	,.R3(R[1676])							,.clk(clk)	,.L(L201)	,.P(P[200])	,.reset(reset)	);
VNU_3 VNU202	(.Q1(Q[122])	,.Q2(Q[584])	,.Q3(Q[1538])							,.R1(R[122])	,.R2(R[584])	,.R3(R[1538])							,.clk(clk)	,.L(L202)	,.P(P[201])	,.reset(reset)	);
VNU_3 VNU203	(.Q1(Q[128])	,.Q2(Q[590])	,.Q3(Q[1544])							,.R1(R[128])	,.R2(R[590])	,.R3(R[1544])							,.clk(clk)	,.L(L203)	,.P(P[202])	,.reset(reset)	);
VNU_3 VNU204	(.Q1(Q[134])	,.Q2(Q[596])	,.Q3(Q[1550])							,.R1(R[134])	,.R2(R[596])	,.R3(R[1550])							,.clk(clk)	,.L(L204)	,.P(P[203])	,.reset(reset)	);
VNU_3 VNU205	(.Q1(Q[140])	,.Q2(Q[602])	,.Q3(Q[1556])							,.R1(R[140])	,.R2(R[602])	,.R3(R[1556])							,.clk(clk)	,.L(L205)	,.P(P[204])	,.reset(reset)	);
VNU_3 VNU206	(.Q1(Q[2])	,.Q2(Q[608])	,.Q3(Q[1562])							,.R1(R[2])	,.R2(R[608])	,.R3(R[1562])							,.clk(clk)	,.L(L206)	,.P(P[205])	,.reset(reset)	);
VNU_3 VNU207	(.Q1(Q[8])	,.Q2(Q[614])	,.Q3(Q[1568])							,.R1(R[8])	,.R2(R[614])	,.R3(R[1568])							,.clk(clk)	,.L(L207)	,.P(P[206])	,.reset(reset)	);
VNU_3 VNU208	(.Q1(Q[14])	,.Q2(Q[620])	,.Q3(Q[1574])							,.R1(R[14])	,.R2(R[620])	,.R3(R[1574])							,.clk(clk)	,.L(L208)	,.P(P[207])	,.reset(reset)	);
VNU_3 VNU209	(.Q1(Q[20])	,.Q2(Q[482])	,.Q3(Q[1580])							,.R1(R[20])	,.R2(R[482])	,.R3(R[1580])							,.clk(clk)	,.L(L209)	,.P(P[208])	,.reset(reset)	);
VNU_3 VNU210	(.Q1(Q[26])	,.Q2(Q[488])	,.Q3(Q[1586])							,.R1(R[26])	,.R2(R[488])	,.R3(R[1586])							,.clk(clk)	,.L(L210)	,.P(P[209])	,.reset(reset)	);
VNU_3 VNU211	(.Q1(Q[32])	,.Q2(Q[494])	,.Q3(Q[1592])							,.R1(R[32])	,.R2(R[494])	,.R3(R[1592])							,.clk(clk)	,.L(L211)	,.P(P[210])	,.reset(reset)	);
VNU_3 VNU212	(.Q1(Q[38])	,.Q2(Q[500])	,.Q3(Q[1598])							,.R1(R[38])	,.R2(R[500])	,.R3(R[1598])							,.clk(clk)	,.L(L212)	,.P(P[211])	,.reset(reset)	);
VNU_3 VNU213	(.Q1(Q[44])	,.Q2(Q[506])	,.Q3(Q[1604])							,.R1(R[44])	,.R2(R[506])	,.R3(R[1604])							,.clk(clk)	,.L(L213)	,.P(P[212])	,.reset(reset)	);
VNU_3 VNU214	(.Q1(Q[50])	,.Q2(Q[512])	,.Q3(Q[1610])							,.R1(R[50])	,.R2(R[512])	,.R3(R[1610])							,.clk(clk)	,.L(L214)	,.P(P[213])	,.reset(reset)	);
VNU_3 VNU215	(.Q1(Q[56])	,.Q2(Q[518])	,.Q3(Q[1616])							,.R1(R[56])	,.R2(R[518])	,.R3(R[1616])							,.clk(clk)	,.L(L215)	,.P(P[214])	,.reset(reset)	);
VNU_3 VNU216	(.Q1(Q[62])	,.Q2(Q[524])	,.Q3(Q[1622])							,.R1(R[62])	,.R2(R[524])	,.R3(R[1622])							,.clk(clk)	,.L(L216)	,.P(P[215])	,.reset(reset)	);
VNU_6 VNU217	(.Q1(Q[27])	,.Q2(Q[591])	,.Q3(Q[710])	,.Q4(Q[1064])	,.Q5(Q[1161])	,.Q6(Q[1611])	,.R1(R[27])	,.R2(R[591])	,.R3(R[710])	,.R4(R[1064])	,.R5(R[1161])	,.R6(R[1611])	,.clk(clk)	,.L(L217)	,.P(P[216])	,.reset(reset)	);
VNU_6 VNU218	(.Q1(Q[33])	,.Q2(Q[597])	,.Q3(Q[716])	,.Q4(Q[1070])	,.Q5(Q[1167])	,.Q6(Q[1617])	,.R1(R[33])	,.R2(R[597])	,.R3(R[716])	,.R4(R[1070])	,.R5(R[1167])	,.R6(R[1617])	,.clk(clk)	,.L(L218)	,.P(P[217])	,.reset(reset)	);
VNU_6 VNU219	(.Q1(Q[39])	,.Q2(Q[603])	,.Q3(Q[722])	,.Q4(Q[1076])	,.Q5(Q[1173])	,.Q6(Q[1623])	,.R1(R[39])	,.R2(R[603])	,.R3(R[722])	,.R4(R[1076])	,.R5(R[1173])	,.R6(R[1623])	,.clk(clk)	,.L(L219)	,.P(P[218])	,.reset(reset)	);
VNU_6 VNU220	(.Q1(Q[45])	,.Q2(Q[609])	,.Q3(Q[728])	,.Q4(Q[938])	,.Q5(Q[1179])	,.Q6(Q[1629])	,.R1(R[45])	,.R2(R[609])	,.R3(R[728])	,.R4(R[938])	,.R5(R[1179])	,.R6(R[1629])	,.clk(clk)	,.L(L220)	,.P(P[219])	,.reset(reset)	);
VNU_6 VNU221	(.Q1(Q[51])	,.Q2(Q[615])	,.Q3(Q[734])	,.Q4(Q[944])	,.Q5(Q[1185])	,.Q6(Q[1635])	,.R1(R[51])	,.R2(R[615])	,.R3(R[734])	,.R4(R[944])	,.R5(R[1185])	,.R6(R[1635])	,.clk(clk)	,.L(L221)	,.P(P[220])	,.reset(reset)	);
VNU_6 VNU222	(.Q1(Q[57])	,.Q2(Q[621])	,.Q3(Q[740])	,.Q4(Q[950])	,.Q5(Q[1191])	,.Q6(Q[1641])	,.R1(R[57])	,.R2(R[621])	,.R3(R[740])	,.R4(R[950])	,.R5(R[1191])	,.R6(R[1641])	,.clk(clk)	,.L(L222)	,.P(P[221])	,.reset(reset)	);
VNU_6 VNU223	(.Q1(Q[63])	,.Q2(Q[483])	,.Q3(Q[746])	,.Q4(Q[956])	,.Q5(Q[1197])	,.Q6(Q[1647])	,.R1(R[63])	,.R2(R[483])	,.R3(R[746])	,.R4(R[956])	,.R5(R[1197])	,.R6(R[1647])	,.clk(clk)	,.L(L223)	,.P(P[222])	,.reset(reset)	);
VNU_6 VNU224	(.Q1(Q[69])	,.Q2(Q[489])	,.Q3(Q[752])	,.Q4(Q[962])	,.Q5(Q[1203])	,.Q6(Q[1653])	,.R1(R[69])	,.R2(R[489])	,.R3(R[752])	,.R4(R[962])	,.R5(R[1203])	,.R6(R[1653])	,.clk(clk)	,.L(L224)	,.P(P[223])	,.reset(reset)	);
VNU_6 VNU225	(.Q1(Q[75])	,.Q2(Q[495])	,.Q3(Q[758])	,.Q4(Q[968])	,.Q5(Q[1209])	,.Q6(Q[1659])	,.R1(R[75])	,.R2(R[495])	,.R3(R[758])	,.R4(R[968])	,.R5(R[1209])	,.R6(R[1659])	,.clk(clk)	,.L(L225)	,.P(P[224])	,.reset(reset)	);
VNU_6 VNU226	(.Q1(Q[81])	,.Q2(Q[501])	,.Q3(Q[764])	,.Q4(Q[974])	,.Q5(Q[1215])	,.Q6(Q[1665])	,.R1(R[81])	,.R2(R[501])	,.R3(R[764])	,.R4(R[974])	,.R5(R[1215])	,.R6(R[1665])	,.clk(clk)	,.L(L226)	,.P(P[225])	,.reset(reset)	);
VNU_6 VNU227	(.Q1(Q[87])	,.Q2(Q[507])	,.Q3(Q[626])	,.Q4(Q[980])	,.Q5(Q[1221])	,.Q6(Q[1671])	,.R1(R[87])	,.R2(R[507])	,.R3(R[626])	,.R4(R[980])	,.R5(R[1221])	,.R6(R[1671])	,.clk(clk)	,.L(L227)	,.P(P[226])	,.reset(reset)	);
VNU_6 VNU228	(.Q1(Q[93])	,.Q2(Q[513])	,.Q3(Q[632])	,.Q4(Q[986])	,.Q5(Q[1083])	,.Q6(Q[1677])	,.R1(R[93])	,.R2(R[513])	,.R3(R[632])	,.R4(R[986])	,.R5(R[1083])	,.R6(R[1677])	,.clk(clk)	,.L(L228)	,.P(P[227])	,.reset(reset)	);
VNU_6 VNU229	(.Q1(Q[99])	,.Q2(Q[519])	,.Q3(Q[638])	,.Q4(Q[992])	,.Q5(Q[1089])	,.Q6(Q[1539])	,.R1(R[99])	,.R2(R[519])	,.R3(R[638])	,.R4(R[992])	,.R5(R[1089])	,.R6(R[1539])	,.clk(clk)	,.L(L229)	,.P(P[228])	,.reset(reset)	);
VNU_6 VNU230	(.Q1(Q[105])	,.Q2(Q[525])	,.Q3(Q[644])	,.Q4(Q[998])	,.Q5(Q[1095])	,.Q6(Q[1545])	,.R1(R[105])	,.R2(R[525])	,.R3(R[644])	,.R4(R[998])	,.R5(R[1095])	,.R6(R[1545])	,.clk(clk)	,.L(L230)	,.P(P[229])	,.reset(reset)	);
VNU_6 VNU231	(.Q1(Q[111])	,.Q2(Q[531])	,.Q3(Q[650])	,.Q4(Q[1004])	,.Q5(Q[1101])	,.Q6(Q[1551])	,.R1(R[111])	,.R2(R[531])	,.R3(R[650])	,.R4(R[1004])	,.R5(R[1101])	,.R6(R[1551])	,.clk(clk)	,.L(L231)	,.P(P[230])	,.reset(reset)	);
VNU_6 VNU232	(.Q1(Q[117])	,.Q2(Q[537])	,.Q3(Q[656])	,.Q4(Q[1010])	,.Q5(Q[1107])	,.Q6(Q[1557])	,.R1(R[117])	,.R2(R[537])	,.R3(R[656])	,.R4(R[1010])	,.R5(R[1107])	,.R6(R[1557])	,.clk(clk)	,.L(L232)	,.P(P[231])	,.reset(reset)	);
VNU_6 VNU233	(.Q1(Q[123])	,.Q2(Q[543])	,.Q3(Q[662])	,.Q4(Q[1016])	,.Q5(Q[1113])	,.Q6(Q[1563])	,.R1(R[123])	,.R2(R[543])	,.R3(R[662])	,.R4(R[1016])	,.R5(R[1113])	,.R6(R[1563])	,.clk(clk)	,.L(L233)	,.P(P[232])	,.reset(reset)	);
VNU_6 VNU234	(.Q1(Q[129])	,.Q2(Q[549])	,.Q3(Q[668])	,.Q4(Q[1022])	,.Q5(Q[1119])	,.Q6(Q[1569])	,.R1(R[129])	,.R2(R[549])	,.R3(R[668])	,.R4(R[1022])	,.R5(R[1119])	,.R6(R[1569])	,.clk(clk)	,.L(L234)	,.P(P[233])	,.reset(reset)	);
VNU_6 VNU235	(.Q1(Q[135])	,.Q2(Q[555])	,.Q3(Q[674])	,.Q4(Q[1028])	,.Q5(Q[1125])	,.Q6(Q[1575])	,.R1(R[135])	,.R2(R[555])	,.R3(R[674])	,.R4(R[1028])	,.R5(R[1125])	,.R6(R[1575])	,.clk(clk)	,.L(L235)	,.P(P[234])	,.reset(reset)	);
VNU_6 VNU236	(.Q1(Q[141])	,.Q2(Q[561])	,.Q3(Q[680])	,.Q4(Q[1034])	,.Q5(Q[1131])	,.Q6(Q[1581])	,.R1(R[141])	,.R2(R[561])	,.R3(R[680])	,.R4(R[1034])	,.R5(R[1131])	,.R6(R[1581])	,.clk(clk)	,.L(L236)	,.P(P[235])	,.reset(reset)	);
VNU_6 VNU237	(.Q1(Q[3])	,.Q2(Q[567])	,.Q3(Q[686])	,.Q4(Q[1040])	,.Q5(Q[1137])	,.Q6(Q[1587])	,.R1(R[3])	,.R2(R[567])	,.R3(R[686])	,.R4(R[1040])	,.R5(R[1137])	,.R6(R[1587])	,.clk(clk)	,.L(L237)	,.P(P[236])	,.reset(reset)	);
VNU_6 VNU238	(.Q1(Q[9])	,.Q2(Q[573])	,.Q3(Q[692])	,.Q4(Q[1046])	,.Q5(Q[1143])	,.Q6(Q[1593])	,.R1(R[9])	,.R2(R[573])	,.R3(R[692])	,.R4(R[1046])	,.R5(R[1143])	,.R6(R[1593])	,.clk(clk)	,.L(L238)	,.P(P[237])	,.reset(reset)	);
VNU_6 VNU239	(.Q1(Q[15])	,.Q2(Q[579])	,.Q3(Q[698])	,.Q4(Q[1052])	,.Q5(Q[1149])	,.Q6(Q[1599])	,.R1(R[15])	,.R2(R[579])	,.R3(R[698])	,.R4(R[1052])	,.R5(R[1149])	,.R6(R[1599])	,.clk(clk)	,.L(L239)	,.P(P[238])	,.reset(reset)	);
VNU_6 VNU240	(.Q1(Q[21])	,.Q2(Q[585])	,.Q3(Q[704])	,.Q4(Q[1058])	,.Q5(Q[1155])	,.Q6(Q[1605])	,.R1(R[21])	,.R2(R[585])	,.R3(R[704])	,.R4(R[1058])	,.R5(R[1155])	,.R6(R[1605])	,.clk(clk)	,.L(L240)	,.P(P[239])	,.reset(reset)	);
VNU_3 VNU241	(.Q1(Q[663])	,.Q2(Q[1059])	,.Q3(Q[1436])							,.R1(R[663])	,.R2(R[1059])	,.R3(R[1436])							,.clk(clk)	,.L(L241)	,.P(P[240])	,.reset(reset)	);
VNU_3 VNU242	(.Q1(Q[669])	,.Q2(Q[1065])	,.Q3(Q[1442])							,.R1(R[669])	,.R2(R[1065])	,.R3(R[1442])							,.clk(clk)	,.L(L242)	,.P(P[241])	,.reset(reset)	);
VNU_3 VNU243	(.Q1(Q[675])	,.Q2(Q[1071])	,.Q3(Q[1448])							,.R1(R[675])	,.R2(R[1071])	,.R3(R[1448])							,.clk(clk)	,.L(L243)	,.P(P[242])	,.reset(reset)	);
VNU_3 VNU244	(.Q1(Q[681])	,.Q2(Q[1077])	,.Q3(Q[1454])							,.R1(R[681])	,.R2(R[1077])	,.R3(R[1454])							,.clk(clk)	,.L(L244)	,.P(P[243])	,.reset(reset)	);
VNU_3 VNU245	(.Q1(Q[687])	,.Q2(Q[939])	,.Q3(Q[1460])							,.R1(R[687])	,.R2(R[939])	,.R3(R[1460])							,.clk(clk)	,.L(L245)	,.P(P[244])	,.reset(reset)	);
VNU_3 VNU246	(.Q1(Q[693])	,.Q2(Q[945])	,.Q3(Q[1466])							,.R1(R[693])	,.R2(R[945])	,.R3(R[1466])							,.clk(clk)	,.L(L246)	,.P(P[245])	,.reset(reset)	);
VNU_3 VNU247	(.Q1(Q[699])	,.Q2(Q[951])	,.Q3(Q[1472])							,.R1(R[699])	,.R2(R[951])	,.R3(R[1472])							,.clk(clk)	,.L(L247)	,.P(P[246])	,.reset(reset)	);
VNU_3 VNU248	(.Q1(Q[705])	,.Q2(Q[957])	,.Q3(Q[1478])							,.R1(R[705])	,.R2(R[957])	,.R3(R[1478])							,.clk(clk)	,.L(L248)	,.P(P[247])	,.reset(reset)	);
VNU_3 VNU249	(.Q1(Q[711])	,.Q2(Q[963])	,.Q3(Q[1484])							,.R1(R[711])	,.R2(R[963])	,.R3(R[1484])							,.clk(clk)	,.L(L249)	,.P(P[248])	,.reset(reset)	);
VNU_3 VNU250	(.Q1(Q[717])	,.Q2(Q[969])	,.Q3(Q[1490])							,.R1(R[717])	,.R2(R[969])	,.R3(R[1490])							,.clk(clk)	,.L(L250)	,.P(P[249])	,.reset(reset)	);
VNU_3 VNU251	(.Q1(Q[723])	,.Q2(Q[975])	,.Q3(Q[1496])							,.R1(R[723])	,.R2(R[975])	,.R3(R[1496])							,.clk(clk)	,.L(L251)	,.P(P[250])	,.reset(reset)	);
VNU_3 VNU252	(.Q1(Q[729])	,.Q2(Q[981])	,.Q3(Q[1502])							,.R1(R[729])	,.R2(R[981])	,.R3(R[1502])							,.clk(clk)	,.L(L252)	,.P(P[251])	,.reset(reset)	);
VNU_3 VNU253	(.Q1(Q[735])	,.Q2(Q[987])	,.Q3(Q[1508])							,.R1(R[735])	,.R2(R[987])	,.R3(R[1508])							,.clk(clk)	,.L(L253)	,.P(P[252])	,.reset(reset)	);
VNU_3 VNU254	(.Q1(Q[741])	,.Q2(Q[993])	,.Q3(Q[1514])							,.R1(R[741])	,.R2(R[993])	,.R3(R[1514])							,.clk(clk)	,.L(L254)	,.P(P[253])	,.reset(reset)	);
VNU_3 VNU255	(.Q1(Q[747])	,.Q2(Q[999])	,.Q3(Q[1520])							,.R1(R[747])	,.R2(R[999])	,.R3(R[1520])							,.clk(clk)	,.L(L255)	,.P(P[254])	,.reset(reset)	);
VNU_3 VNU256	(.Q1(Q[753])	,.Q2(Q[1005])	,.Q3(Q[1526])							,.R1(R[753])	,.R2(R[1005])	,.R3(R[1526])							,.clk(clk)	,.L(L256)	,.P(P[255])	,.reset(reset)	);
VNU_3 VNU257	(.Q1(Q[759])	,.Q2(Q[1011])	,.Q3(Q[1532])							,.R1(R[759])	,.R2(R[1011])	,.R3(R[1532])							,.clk(clk)	,.L(L257)	,.P(P[256])	,.reset(reset)	);
VNU_3 VNU258	(.Q1(Q[765])	,.Q2(Q[1017])	,.Q3(Q[1394])							,.R1(R[765])	,.R2(R[1017])	,.R3(R[1394])							,.clk(clk)	,.L(L258)	,.P(P[257])	,.reset(reset)	);
VNU_3 VNU259	(.Q1(Q[627])	,.Q2(Q[1023])	,.Q3(Q[1400])							,.R1(R[627])	,.R2(R[1023])	,.R3(R[1400])							,.clk(clk)	,.L(L259)	,.P(P[258])	,.reset(reset)	);
VNU_3 VNU260	(.Q1(Q[633])	,.Q2(Q[1029])	,.Q3(Q[1406])							,.R1(R[633])	,.R2(R[1029])	,.R3(R[1406])							,.clk(clk)	,.L(L260)	,.P(P[259])	,.reset(reset)	);
VNU_3 VNU261	(.Q1(Q[639])	,.Q2(Q[1035])	,.Q3(Q[1412])							,.R1(R[639])	,.R2(R[1035])	,.R3(R[1412])							,.clk(clk)	,.L(L261)	,.P(P[260])	,.reset(reset)	);
VNU_3 VNU262	(.Q1(Q[645])	,.Q2(Q[1041])	,.Q3(Q[1418])							,.R1(R[645])	,.R2(R[1041])	,.R3(R[1418])							,.clk(clk)	,.L(L262)	,.P(P[261])	,.reset(reset)	);
VNU_3 VNU263	(.Q1(Q[651])	,.Q2(Q[1047])	,.Q3(Q[1424])							,.R1(R[651])	,.R2(R[1047])	,.R3(R[1424])							,.clk(clk)	,.L(L263)	,.P(P[262])	,.reset(reset)	);
VNU_3 VNU264	(.Q1(Q[657])	,.Q2(Q[1053])	,.Q3(Q[1430])							,.R1(R[657])	,.R2(R[1053])	,.R3(R[1430])							,.clk(clk)	,.L(L264)	,.P(P[263])	,.reset(reset)	);
VNU_6 VNU265	(.Q1(Q[295])	,.Q2(Q[316])	,.Q3(Q[806])	,.Q4(Q[1312])	,.Q5(Q[1431])	,.Q6(Q[1791])	,.R1(R[295])	,.R2(R[316])	,.R3(R[806])	,.R4(R[1312])	,.R5(R[1431])	,.R6(R[1791])	,.clk(clk)	,.L(L265)	,.P(P[264])	,.reset(reset)	);
VNU_6 VNU266	(.Q1(Q[302])	,.Q2(Q[323])	,.Q3(Q[813])	,.Q4(Q[1319])	,.Q5(Q[1437])	,.Q6(Q[1797])	,.R1(R[302])	,.R2(R[323])	,.R3(R[813])	,.R4(R[1319])	,.R5(R[1437])	,.R6(R[1797])	,.clk(clk)	,.L(L266)	,.P(P[265])	,.reset(reset)	);
VNU_6 VNU267	(.Q1(Q[309])	,.Q2(Q[330])	,.Q3(Q[820])	,.Q4(Q[1326])	,.Q5(Q[1443])	,.Q6(Q[1803])	,.R1(R[309])	,.R2(R[330])	,.R3(R[820])	,.R4(R[1326])	,.R5(R[1443])	,.R6(R[1803])	,.clk(clk)	,.L(L267)	,.P(P[266])	,.reset(reset)	);
VNU_6 VNU268	(.Q1(Q[148])	,.Q2(Q[337])	,.Q3(Q[827])	,.Q4(Q[1333])	,.Q5(Q[1449])	,.Q6(Q[1809])	,.R1(R[148])	,.R2(R[337])	,.R3(R[827])	,.R4(R[1333])	,.R5(R[1449])	,.R6(R[1809])	,.clk(clk)	,.L(L268)	,.P(P[267])	,.reset(reset)	);
VNU_6 VNU269	(.Q1(Q[155])	,.Q2(Q[344])	,.Q3(Q[834])	,.Q4(Q[1340])	,.Q5(Q[1455])	,.Q6(Q[1815])	,.R1(R[155])	,.R2(R[344])	,.R3(R[834])	,.R4(R[1340])	,.R5(R[1455])	,.R6(R[1815])	,.clk(clk)	,.L(L269)	,.P(P[268])	,.reset(reset)	);
VNU_6 VNU270	(.Q1(Q[162])	,.Q2(Q[351])	,.Q3(Q[841])	,.Q4(Q[1347])	,.Q5(Q[1461])	,.Q6(Q[1821])	,.R1(R[162])	,.R2(R[351])	,.R3(R[841])	,.R4(R[1347])	,.R5(R[1461])	,.R6(R[1821])	,.clk(clk)	,.L(L270)	,.P(P[269])	,.reset(reset)	);
VNU_6 VNU271	(.Q1(Q[169])	,.Q2(Q[358])	,.Q3(Q[848])	,.Q4(Q[1354])	,.Q5(Q[1467])	,.Q6(Q[1683])	,.R1(R[169])	,.R2(R[358])	,.R3(R[848])	,.R4(R[1354])	,.R5(R[1467])	,.R6(R[1683])	,.clk(clk)	,.L(L271)	,.P(P[270])	,.reset(reset)	);
VNU_6 VNU272	(.Q1(Q[176])	,.Q2(Q[365])	,.Q3(Q[855])	,.Q4(Q[1361])	,.Q5(Q[1473])	,.Q6(Q[1689])	,.R1(R[176])	,.R2(R[365])	,.R3(R[855])	,.R4(R[1361])	,.R5(R[1473])	,.R6(R[1689])	,.clk(clk)	,.L(L272)	,.P(P[271])	,.reset(reset)	);
VNU_6 VNU273	(.Q1(Q[183])	,.Q2(Q[372])	,.Q3(Q[862])	,.Q4(Q[1368])	,.Q5(Q[1479])	,.Q6(Q[1695])	,.R1(R[183])	,.R2(R[372])	,.R3(R[862])	,.R4(R[1368])	,.R5(R[1479])	,.R6(R[1695])	,.clk(clk)	,.L(L273)	,.P(P[272])	,.reset(reset)	);
VNU_6 VNU274	(.Q1(Q[190])	,.Q2(Q[379])	,.Q3(Q[869])	,.Q4(Q[1375])	,.Q5(Q[1485])	,.Q6(Q[1701])	,.R1(R[190])	,.R2(R[379])	,.R3(R[869])	,.R4(R[1375])	,.R5(R[1485])	,.R6(R[1701])	,.clk(clk)	,.L(L274)	,.P(P[273])	,.reset(reset)	);
VNU_6 VNU275	(.Q1(Q[197])	,.Q2(Q[386])	,.Q3(Q[876])	,.Q4(Q[1382])	,.Q5(Q[1491])	,.Q6(Q[1707])	,.R1(R[197])	,.R2(R[386])	,.R3(R[876])	,.R4(R[1382])	,.R5(R[1491])	,.R6(R[1707])	,.clk(clk)	,.L(L275)	,.P(P[274])	,.reset(reset)	);
VNU_6 VNU276	(.Q1(Q[204])	,.Q2(Q[393])	,.Q3(Q[883])	,.Q4(Q[1389])	,.Q5(Q[1497])	,.Q6(Q[1713])	,.R1(R[204])	,.R2(R[393])	,.R3(R[883])	,.R4(R[1389])	,.R5(R[1497])	,.R6(R[1713])	,.clk(clk)	,.L(L276)	,.P(P[275])	,.reset(reset)	);
VNU_6 VNU277	(.Q1(Q[211])	,.Q2(Q[400])	,.Q3(Q[890])	,.Q4(Q[1228])	,.Q5(Q[1503])	,.Q6(Q[1719])	,.R1(R[211])	,.R2(R[400])	,.R3(R[890])	,.R4(R[1228])	,.R5(R[1503])	,.R6(R[1719])	,.clk(clk)	,.L(L277)	,.P(P[276])	,.reset(reset)	);
VNU_6 VNU278	(.Q1(Q[218])	,.Q2(Q[407])	,.Q3(Q[897])	,.Q4(Q[1235])	,.Q5(Q[1509])	,.Q6(Q[1725])	,.R1(R[218])	,.R2(R[407])	,.R3(R[897])	,.R4(R[1235])	,.R5(R[1509])	,.R6(R[1725])	,.clk(clk)	,.L(L278)	,.P(P[277])	,.reset(reset)	);
VNU_6 VNU279	(.Q1(Q[225])	,.Q2(Q[414])	,.Q3(Q[904])	,.Q4(Q[1242])	,.Q5(Q[1515])	,.Q6(Q[1731])	,.R1(R[225])	,.R2(R[414])	,.R3(R[904])	,.R4(R[1242])	,.R5(R[1515])	,.R6(R[1731])	,.clk(clk)	,.L(L279)	,.P(P[278])	,.reset(reset)	);
VNU_6 VNU280	(.Q1(Q[232])	,.Q2(Q[421])	,.Q3(Q[911])	,.Q4(Q[1249])	,.Q5(Q[1521])	,.Q6(Q[1737])	,.R1(R[232])	,.R2(R[421])	,.R3(R[911])	,.R4(R[1249])	,.R5(R[1521])	,.R6(R[1737])	,.clk(clk)	,.L(L280)	,.P(P[279])	,.reset(reset)	);
VNU_6 VNU281	(.Q1(Q[239])	,.Q2(Q[428])	,.Q3(Q[918])	,.Q4(Q[1256])	,.Q5(Q[1527])	,.Q6(Q[1743])	,.R1(R[239])	,.R2(R[428])	,.R3(R[918])	,.R4(R[1256])	,.R5(R[1527])	,.R6(R[1743])	,.clk(clk)	,.L(L281)	,.P(P[280])	,.reset(reset)	);
VNU_6 VNU282	(.Q1(Q[246])	,.Q2(Q[435])	,.Q3(Q[925])	,.Q4(Q[1263])	,.Q5(Q[1533])	,.Q6(Q[1749])	,.R1(R[246])	,.R2(R[435])	,.R3(R[925])	,.R4(R[1263])	,.R5(R[1533])	,.R6(R[1749])	,.clk(clk)	,.L(L282)	,.P(P[281])	,.reset(reset)	);
VNU_6 VNU283	(.Q1(Q[253])	,.Q2(Q[442])	,.Q3(Q[932])	,.Q4(Q[1270])	,.Q5(Q[1395])	,.Q6(Q[1755])	,.R1(R[253])	,.R2(R[442])	,.R3(R[932])	,.R4(R[1270])	,.R5(R[1395])	,.R6(R[1755])	,.clk(clk)	,.L(L283)	,.P(P[282])	,.reset(reset)	);
VNU_6 VNU284	(.Q1(Q[260])	,.Q2(Q[449])	,.Q3(Q[771])	,.Q4(Q[1277])	,.Q5(Q[1401])	,.Q6(Q[1761])	,.R1(R[260])	,.R2(R[449])	,.R3(R[771])	,.R4(R[1277])	,.R5(R[1401])	,.R6(R[1761])	,.clk(clk)	,.L(L284)	,.P(P[283])	,.reset(reset)	);
VNU_6 VNU285	(.Q1(Q[267])	,.Q2(Q[456])	,.Q3(Q[778])	,.Q4(Q[1284])	,.Q5(Q[1407])	,.Q6(Q[1767])	,.R1(R[267])	,.R2(R[456])	,.R3(R[778])	,.R4(R[1284])	,.R5(R[1407])	,.R6(R[1767])	,.clk(clk)	,.L(L285)	,.P(P[284])	,.reset(reset)	);
VNU_6 VNU286	(.Q1(Q[274])	,.Q2(Q[463])	,.Q3(Q[785])	,.Q4(Q[1291])	,.Q5(Q[1413])	,.Q6(Q[1773])	,.R1(R[274])	,.R2(R[463])	,.R3(R[785])	,.R4(R[1291])	,.R5(R[1413])	,.R6(R[1773])	,.clk(clk)	,.L(L286)	,.P(P[285])	,.reset(reset)	);
VNU_6 VNU287	(.Q1(Q[281])	,.Q2(Q[470])	,.Q3(Q[792])	,.Q4(Q[1298])	,.Q5(Q[1419])	,.Q6(Q[1779])	,.R1(R[281])	,.R2(R[470])	,.R3(R[792])	,.R4(R[1298])	,.R5(R[1419])	,.R6(R[1779])	,.clk(clk)	,.L(L287)	,.P(P[286])	,.reset(reset)	);
VNU_6 VNU288	(.Q1(Q[288])	,.Q2(Q[477])	,.Q3(Q[799])	,.Q4(Q[1305])	,.Q5(Q[1425])	,.Q6(Q[1785])	,.R1(R[288])	,.R2(R[477])	,.R3(R[799])	,.R4(R[1305])	,.R5(R[1425])	,.R6(R[1785])	,.clk(clk)	,.L(L288)	,.P(P[287])	,.reset(reset)	);
VNU_3 VNU289	(.Q1(Q[142])	,.Q2(Q[772])	,.Q3(Q[1822])							,.R1(R[142])	,.R2(R[772])	,.R3(R[1822])							,.clk(clk)	,.L(L289)	,.P(P[288])	,.reset(reset)	);
VNU_3 VNU290	(.Q1(Q[4])	,.Q2(Q[779])	,.Q3(Q[1684])							,.R1(R[4])	,.R2(R[779])	,.R3(R[1684])							,.clk(clk)	,.L(L290)	,.P(P[289])	,.reset(reset)	);
VNU_3 VNU291	(.Q1(Q[10])	,.Q2(Q[786])	,.Q3(Q[1690])							,.R1(R[10])	,.R2(R[786])	,.R3(R[1690])							,.clk(clk)	,.L(L291)	,.P(P[290])	,.reset(reset)	);
VNU_3 VNU292	(.Q1(Q[16])	,.Q2(Q[793])	,.Q3(Q[1696])							,.R1(R[16])	,.R2(R[793])	,.R3(R[1696])							,.clk(clk)	,.L(L292)	,.P(P[291])	,.reset(reset)	);
VNU_3 VNU293	(.Q1(Q[22])	,.Q2(Q[800])	,.Q3(Q[1702])							,.R1(R[22])	,.R2(R[800])	,.R3(R[1702])							,.clk(clk)	,.L(L293)	,.P(P[292])	,.reset(reset)	);
VNU_3 VNU294	(.Q1(Q[28])	,.Q2(Q[807])	,.Q3(Q[1708])							,.R1(R[28])	,.R2(R[807])	,.R3(R[1708])							,.clk(clk)	,.L(L294)	,.P(P[293])	,.reset(reset)	);
VNU_3 VNU295	(.Q1(Q[34])	,.Q2(Q[814])	,.Q3(Q[1714])							,.R1(R[34])	,.R2(R[814])	,.R3(R[1714])							,.clk(clk)	,.L(L295)	,.P(P[294])	,.reset(reset)	);
VNU_3 VNU296	(.Q1(Q[40])	,.Q2(Q[821])	,.Q3(Q[1720])							,.R1(R[40])	,.R2(R[821])	,.R3(R[1720])							,.clk(clk)	,.L(L296)	,.P(P[295])	,.reset(reset)	);
VNU_3 VNU297	(.Q1(Q[46])	,.Q2(Q[828])	,.Q3(Q[1726])							,.R1(R[46])	,.R2(R[828])	,.R3(R[1726])							,.clk(clk)	,.L(L297)	,.P(P[296])	,.reset(reset)	);
VNU_3 VNU298	(.Q1(Q[52])	,.Q2(Q[835])	,.Q3(Q[1732])							,.R1(R[52])	,.R2(R[835])	,.R3(R[1732])							,.clk(clk)	,.L(L298)	,.P(P[297])	,.reset(reset)	);
VNU_3 VNU299	(.Q1(Q[58])	,.Q2(Q[842])	,.Q3(Q[1738])							,.R1(R[58])	,.R2(R[842])	,.R3(R[1738])							,.clk(clk)	,.L(L299)	,.P(P[298])	,.reset(reset)	);
VNU_3 VNU300	(.Q1(Q[64])	,.Q2(Q[849])	,.Q3(Q[1744])							,.R1(R[64])	,.R2(R[849])	,.R3(R[1744])							,.clk(clk)	,.L(L300)	,.P(P[299])	,.reset(reset)	);
VNU_3 VNU301	(.Q1(Q[70])	,.Q2(Q[856])	,.Q3(Q[1750])							,.R1(R[70])	,.R2(R[856])	,.R3(R[1750])							,.clk(clk)	,.L(L301)	,.P(P[300])	,.reset(reset)	);
VNU_3 VNU302	(.Q1(Q[76])	,.Q2(Q[863])	,.Q3(Q[1756])							,.R1(R[76])	,.R2(R[863])	,.R3(R[1756])							,.clk(clk)	,.L(L302)	,.P(P[301])	,.reset(reset)	);
VNU_3 VNU303	(.Q1(Q[82])	,.Q2(Q[870])	,.Q3(Q[1762])							,.R1(R[82])	,.R2(R[870])	,.R3(R[1762])							,.clk(clk)	,.L(L303)	,.P(P[302])	,.reset(reset)	);
VNU_3 VNU304	(.Q1(Q[88])	,.Q2(Q[877])	,.Q3(Q[1768])							,.R1(R[88])	,.R2(R[877])	,.R3(R[1768])							,.clk(clk)	,.L(L304)	,.P(P[303])	,.reset(reset)	);
VNU_3 VNU305	(.Q1(Q[94])	,.Q2(Q[884])	,.Q3(Q[1774])							,.R1(R[94])	,.R2(R[884])	,.R3(R[1774])							,.clk(clk)	,.L(L305)	,.P(P[304])	,.reset(reset)	);
VNU_3 VNU306	(.Q1(Q[100])	,.Q2(Q[891])	,.Q3(Q[1780])							,.R1(R[100])	,.R2(R[891])	,.R3(R[1780])							,.clk(clk)	,.L(L306)	,.P(P[305])	,.reset(reset)	);
VNU_3 VNU307	(.Q1(Q[106])	,.Q2(Q[898])	,.Q3(Q[1786])							,.R1(R[106])	,.R2(R[898])	,.R3(R[1786])							,.clk(clk)	,.L(L307)	,.P(P[306])	,.reset(reset)	);
VNU_3 VNU308	(.Q1(Q[112])	,.Q2(Q[905])	,.Q3(Q[1792])							,.R1(R[112])	,.R2(R[905])	,.R3(R[1792])							,.clk(clk)	,.L(L308)	,.P(P[307])	,.reset(reset)	);
VNU_3 VNU309	(.Q1(Q[118])	,.Q2(Q[912])	,.Q3(Q[1798])							,.R1(R[118])	,.R2(R[912])	,.R3(R[1798])							,.clk(clk)	,.L(L309)	,.P(P[308])	,.reset(reset)	);
VNU_3 VNU310	(.Q1(Q[124])	,.Q2(Q[919])	,.Q3(Q[1804])							,.R1(R[124])	,.R2(R[919])	,.R3(R[1804])							,.clk(clk)	,.L(L310)	,.P(P[309])	,.reset(reset)	);
VNU_3 VNU311	(.Q1(Q[130])	,.Q2(Q[926])	,.Q3(Q[1810])							,.R1(R[130])	,.R2(R[926])	,.R3(R[1810])							,.clk(clk)	,.L(L311)	,.P(P[310])	,.reset(reset)	);
VNU_3 VNU312	(.Q1(Q[136])	,.Q2(Q[933])	,.Q3(Q[1816])							,.R1(R[136])	,.R2(R[933])	,.R3(R[1816])							,.clk(clk)	,.L(L312)	,.P(P[311])	,.reset(reset)	);
VNU_2 VNU313	(.Q1(Q[5])	,.Q2(Q[149])									,.R1(R[5])	,.R2(R[149])									,.clk(clk)	,.L(L313)	,.P(P[312])	,.reset(reset)	);
VNU_2 VNU314	(.Q1(Q[11])	,.Q2(Q[156])									,.R1(R[11])	,.R2(R[156])									,.clk(clk)	,.L(L314)	,.P(P[313])	,.reset(reset)	);
VNU_2 VNU315	(.Q1(Q[17])	,.Q2(Q[163])									,.R1(R[17])	,.R2(R[163])									,.clk(clk)	,.L(L315)	,.P(P[314])	,.reset(reset)	);
VNU_2 VNU316	(.Q1(Q[23])	,.Q2(Q[170])									,.R1(R[23])	,.R2(R[170])									,.clk(clk)	,.L(L316)	,.P(P[315])	,.reset(reset)	);
VNU_2 VNU317	(.Q1(Q[29])	,.Q2(Q[177])									,.R1(R[29])	,.R2(R[177])									,.clk(clk)	,.L(L317)	,.P(P[316])	,.reset(reset)	);
VNU_2 VNU318	(.Q1(Q[35])	,.Q2(Q[184])									,.R1(R[35])	,.R2(R[184])									,.clk(clk)	,.L(L318)	,.P(P[317])	,.reset(reset)	);
VNU_2 VNU319	(.Q1(Q[41])	,.Q2(Q[191])									,.R1(R[41])	,.R2(R[191])									,.clk(clk)	,.L(L319)	,.P(P[318])	,.reset(reset)	);
VNU_2 VNU320	(.Q1(Q[47])	,.Q2(Q[198])									,.R1(R[47])	,.R2(R[198])									,.clk(clk)	,.L(L320)	,.P(P[319])	,.reset(reset)	);
VNU_2 VNU321	(.Q1(Q[53])	,.Q2(Q[205])									,.R1(R[53])	,.R2(R[205])									,.clk(clk)	,.L(L321)	,.P(P[320])	,.reset(reset)	);
VNU_2 VNU322	(.Q1(Q[59])	,.Q2(Q[212])									,.R1(R[59])	,.R2(R[212])									,.clk(clk)	,.L(L322)	,.P(P[321])	,.reset(reset)	);
VNU_2 VNU323	(.Q1(Q[65])	,.Q2(Q[219])									,.R1(R[65])	,.R2(R[219])									,.clk(clk)	,.L(L323)	,.P(P[322])	,.reset(reset)	);
VNU_2 VNU324	(.Q1(Q[71])	,.Q2(Q[226])									,.R1(R[71])	,.R2(R[226])									,.clk(clk)	,.L(L324)	,.P(P[323])	,.reset(reset)	);
VNU_2 VNU325	(.Q1(Q[77])	,.Q2(Q[233])									,.R1(R[77])	,.R2(R[233])									,.clk(clk)	,.L(L325)	,.P(P[324])	,.reset(reset)	);
VNU_2 VNU326	(.Q1(Q[83])	,.Q2(Q[240])									,.R1(R[83])	,.R2(R[240])									,.clk(clk)	,.L(L326)	,.P(P[325])	,.reset(reset)	);
VNU_2 VNU327	(.Q1(Q[89])	,.Q2(Q[247])									,.R1(R[89])	,.R2(R[247])									,.clk(clk)	,.L(L327)	,.P(P[326])	,.reset(reset)	);
VNU_2 VNU328	(.Q1(Q[95])	,.Q2(Q[254])									,.R1(R[95])	,.R2(R[254])									,.clk(clk)	,.L(L328)	,.P(P[327])	,.reset(reset)	);
VNU_2 VNU329	(.Q1(Q[101])	,.Q2(Q[261])									,.R1(R[101])	,.R2(R[261])									,.clk(clk)	,.L(L329)	,.P(P[328])	,.reset(reset)	);
VNU_2 VNU330	(.Q1(Q[107])	,.Q2(Q[268])									,.R1(R[107])	,.R2(R[268])									,.clk(clk)	,.L(L330)	,.P(P[329])	,.reset(reset)	);
VNU_2 VNU331	(.Q1(Q[113])	,.Q2(Q[275])									,.R1(R[113])	,.R2(R[275])									,.clk(clk)	,.L(L331)	,.P(P[330])	,.reset(reset)	);
VNU_2 VNU332	(.Q1(Q[119])	,.Q2(Q[282])									,.R1(R[119])	,.R2(R[282])									,.clk(clk)	,.L(L332)	,.P(P[331])	,.reset(reset)	);
VNU_2 VNU333	(.Q1(Q[125])	,.Q2(Q[289])									,.R1(R[125])	,.R2(R[289])									,.clk(clk)	,.L(L333)	,.P(P[332])	,.reset(reset)	);
VNU_2 VNU334	(.Q1(Q[131])	,.Q2(Q[296])									,.R1(R[131])	,.R2(R[296])									,.clk(clk)	,.L(L334)	,.P(P[333])	,.reset(reset)	);
VNU_2 VNU335	(.Q1(Q[137])	,.Q2(Q[303])									,.R1(R[137])	,.R2(R[303])									,.clk(clk)	,.L(L335)	,.P(P[334])	,.reset(reset)	);
VNU_2 VNU336	(.Q1(Q[143])	,.Q2(Q[310])									,.R1(R[143])	,.R2(R[310])									,.clk(clk)	,.L(L336)	,.P(P[335])	,.reset(reset)	);
VNU_2 VNU337	(.Q1(Q[150])	,.Q2(Q[317])									,.R1(R[150])	,.R2(R[317])									,.clk(clk)	,.L(L337)	,.P(P[336])	,.reset(reset)	);
VNU_2 VNU338	(.Q1(Q[157])	,.Q2(Q[324])									,.R1(R[157])	,.R2(R[324])									,.clk(clk)	,.L(L338)	,.P(P[337])	,.reset(reset)	);
VNU_2 VNU339	(.Q1(Q[164])	,.Q2(Q[331])									,.R1(R[164])	,.R2(R[331])									,.clk(clk)	,.L(L339)	,.P(P[338])	,.reset(reset)	);
VNU_2 VNU340	(.Q1(Q[171])	,.Q2(Q[338])									,.R1(R[171])	,.R2(R[338])									,.clk(clk)	,.L(L340)	,.P(P[339])	,.reset(reset)	);
VNU_2 VNU341	(.Q1(Q[178])	,.Q2(Q[345])									,.R1(R[178])	,.R2(R[345])									,.clk(clk)	,.L(L341)	,.P(P[340])	,.reset(reset)	);
VNU_2 VNU342	(.Q1(Q[185])	,.Q2(Q[352])									,.R1(R[185])	,.R2(R[352])									,.clk(clk)	,.L(L342)	,.P(P[341])	,.reset(reset)	);
VNU_2 VNU343	(.Q1(Q[192])	,.Q2(Q[359])									,.R1(R[192])	,.R2(R[359])									,.clk(clk)	,.L(L343)	,.P(P[342])	,.reset(reset)	);
VNU_2 VNU344	(.Q1(Q[199])	,.Q2(Q[366])									,.R1(R[199])	,.R2(R[366])									,.clk(clk)	,.L(L344)	,.P(P[343])	,.reset(reset)	);
VNU_2 VNU345	(.Q1(Q[206])	,.Q2(Q[373])									,.R1(R[206])	,.R2(R[373])									,.clk(clk)	,.L(L345)	,.P(P[344])	,.reset(reset)	);
VNU_2 VNU346	(.Q1(Q[213])	,.Q2(Q[380])									,.R1(R[213])	,.R2(R[380])									,.clk(clk)	,.L(L346)	,.P(P[345])	,.reset(reset)	);
VNU_2 VNU347	(.Q1(Q[220])	,.Q2(Q[387])									,.R1(R[220])	,.R2(R[387])									,.clk(clk)	,.L(L347)	,.P(P[346])	,.reset(reset)	);
VNU_2 VNU348	(.Q1(Q[227])	,.Q2(Q[394])									,.R1(R[227])	,.R2(R[394])									,.clk(clk)	,.L(L348)	,.P(P[347])	,.reset(reset)	);
VNU_2 VNU349	(.Q1(Q[234])	,.Q2(Q[401])									,.R1(R[234])	,.R2(R[401])									,.clk(clk)	,.L(L349)	,.P(P[348])	,.reset(reset)	);
VNU_2 VNU350	(.Q1(Q[241])	,.Q2(Q[408])									,.R1(R[241])	,.R2(R[408])									,.clk(clk)	,.L(L350)	,.P(P[349])	,.reset(reset)	);
VNU_2 VNU351	(.Q1(Q[248])	,.Q2(Q[415])									,.R1(R[248])	,.R2(R[415])									,.clk(clk)	,.L(L351)	,.P(P[350])	,.reset(reset)	);
VNU_2 VNU352	(.Q1(Q[255])	,.Q2(Q[422])									,.R1(R[255])	,.R2(R[422])									,.clk(clk)	,.L(L352)	,.P(P[351])	,.reset(reset)	);
VNU_2 VNU353	(.Q1(Q[262])	,.Q2(Q[429])									,.R1(R[262])	,.R2(R[429])									,.clk(clk)	,.L(L353)	,.P(P[352])	,.reset(reset)	);
VNU_2 VNU354	(.Q1(Q[269])	,.Q2(Q[436])									,.R1(R[269])	,.R2(R[436])									,.clk(clk)	,.L(L354)	,.P(P[353])	,.reset(reset)	);
VNU_2 VNU355	(.Q1(Q[276])	,.Q2(Q[443])									,.R1(R[276])	,.R2(R[443])									,.clk(clk)	,.L(L355)	,.P(P[354])	,.reset(reset)	);
VNU_2 VNU356	(.Q1(Q[283])	,.Q2(Q[450])									,.R1(R[283])	,.R2(R[450])									,.clk(clk)	,.L(L356)	,.P(P[355])	,.reset(reset)	);
VNU_2 VNU357	(.Q1(Q[290])	,.Q2(Q[457])									,.R1(R[290])	,.R2(R[457])									,.clk(clk)	,.L(L357)	,.P(P[356])	,.reset(reset)	);
VNU_2 VNU358	(.Q1(Q[297])	,.Q2(Q[464])									,.R1(R[297])	,.R2(R[464])									,.clk(clk)	,.L(L358)	,.P(P[357])	,.reset(reset)	);
VNU_2 VNU359	(.Q1(Q[304])	,.Q2(Q[471])									,.R1(R[304])	,.R2(R[471])									,.clk(clk)	,.L(L359)	,.P(P[358])	,.reset(reset)	);
VNU_2 VNU360	(.Q1(Q[311])	,.Q2(Q[478])									,.R1(R[311])	,.R2(R[478])									,.clk(clk)	,.L(L360)	,.P(P[359])	,.reset(reset)	);
VNU_2 VNU361	(.Q1(Q[318])	,.Q2(Q[484])									,.R1(R[318])	,.R2(R[484])									,.clk(clk)	,.L(L361)	,.P(P[360])	,.reset(reset)	);
VNU_2 VNU362	(.Q1(Q[325])	,.Q2(Q[490])									,.R1(R[325])	,.R2(R[490])									,.clk(clk)	,.L(L362)	,.P(P[361])	,.reset(reset)	);
VNU_2 VNU363	(.Q1(Q[332])	,.Q2(Q[496])									,.R1(R[332])	,.R2(R[496])									,.clk(clk)	,.L(L363)	,.P(P[362])	,.reset(reset)	);
VNU_2 VNU364	(.Q1(Q[339])	,.Q2(Q[502])									,.R1(R[339])	,.R2(R[502])									,.clk(clk)	,.L(L364)	,.P(P[363])	,.reset(reset)	);
VNU_2 VNU365	(.Q1(Q[346])	,.Q2(Q[508])									,.R1(R[346])	,.R2(R[508])									,.clk(clk)	,.L(L365)	,.P(P[364])	,.reset(reset)	);
VNU_2 VNU366	(.Q1(Q[353])	,.Q2(Q[514])									,.R1(R[353])	,.R2(R[514])									,.clk(clk)	,.L(L366)	,.P(P[365])	,.reset(reset)	);
VNU_2 VNU367	(.Q1(Q[360])	,.Q2(Q[520])									,.R1(R[360])	,.R2(R[520])									,.clk(clk)	,.L(L367)	,.P(P[366])	,.reset(reset)	);
VNU_2 VNU368	(.Q1(Q[367])	,.Q2(Q[526])									,.R1(R[367])	,.R2(R[526])									,.clk(clk)	,.L(L368)	,.P(P[367])	,.reset(reset)	);
VNU_2 VNU369	(.Q1(Q[374])	,.Q2(Q[532])									,.R1(R[374])	,.R2(R[532])									,.clk(clk)	,.L(L369)	,.P(P[368])	,.reset(reset)	);
VNU_2 VNU370	(.Q1(Q[381])	,.Q2(Q[538])									,.R1(R[381])	,.R2(R[538])									,.clk(clk)	,.L(L370)	,.P(P[369])	,.reset(reset)	);
VNU_2 VNU371	(.Q1(Q[388])	,.Q2(Q[544])									,.R1(R[388])	,.R2(R[544])									,.clk(clk)	,.L(L371)	,.P(P[370])	,.reset(reset)	);
VNU_2 VNU372	(.Q1(Q[395])	,.Q2(Q[550])									,.R1(R[395])	,.R2(R[550])									,.clk(clk)	,.L(L372)	,.P(P[371])	,.reset(reset)	);
VNU_2 VNU373	(.Q1(Q[402])	,.Q2(Q[556])									,.R1(R[402])	,.R2(R[556])									,.clk(clk)	,.L(L373)	,.P(P[372])	,.reset(reset)	);
VNU_2 VNU374	(.Q1(Q[409])	,.Q2(Q[562])									,.R1(R[409])	,.R2(R[562])									,.clk(clk)	,.L(L374)	,.P(P[373])	,.reset(reset)	);
VNU_2 VNU375	(.Q1(Q[416])	,.Q2(Q[568])									,.R1(R[416])	,.R2(R[568])									,.clk(clk)	,.L(L375)	,.P(P[374])	,.reset(reset)	);
VNU_2 VNU376	(.Q1(Q[423])	,.Q2(Q[574])									,.R1(R[423])	,.R2(R[574])									,.clk(clk)	,.L(L376)	,.P(P[375])	,.reset(reset)	);
VNU_2 VNU377	(.Q1(Q[430])	,.Q2(Q[580])									,.R1(R[430])	,.R2(R[580])									,.clk(clk)	,.L(L377)	,.P(P[376])	,.reset(reset)	);
VNU_2 VNU378	(.Q1(Q[437])	,.Q2(Q[586])									,.R1(R[437])	,.R2(R[586])									,.clk(clk)	,.L(L378)	,.P(P[377])	,.reset(reset)	);
VNU_2 VNU379	(.Q1(Q[444])	,.Q2(Q[592])									,.R1(R[444])	,.R2(R[592])									,.clk(clk)	,.L(L379)	,.P(P[378])	,.reset(reset)	);
VNU_2 VNU380	(.Q1(Q[451])	,.Q2(Q[598])									,.R1(R[451])	,.R2(R[598])									,.clk(clk)	,.L(L380)	,.P(P[379])	,.reset(reset)	);
VNU_2 VNU381	(.Q1(Q[458])	,.Q2(Q[604])									,.R1(R[458])	,.R2(R[604])									,.clk(clk)	,.L(L381)	,.P(P[380])	,.reset(reset)	);
VNU_2 VNU382	(.Q1(Q[465])	,.Q2(Q[610])									,.R1(R[465])	,.R2(R[610])									,.clk(clk)	,.L(L382)	,.P(P[381])	,.reset(reset)	);
VNU_2 VNU383	(.Q1(Q[472])	,.Q2(Q[616])									,.R1(R[472])	,.R2(R[616])									,.clk(clk)	,.L(L383)	,.P(P[382])	,.reset(reset)	);
VNU_2 VNU384	(.Q1(Q[479])	,.Q2(Q[622])									,.R1(R[479])	,.R2(R[622])									,.clk(clk)	,.L(L384)	,.P(P[383])	,.reset(reset)	);
VNU_2 VNU385	(.Q1(Q[485])	,.Q2(Q[628])									,.R1(R[485])	,.R2(R[628])									,.clk(clk)	,.L(L385)	,.P(P[384])	,.reset(reset)	);
VNU_2 VNU386	(.Q1(Q[491])	,.Q2(Q[634])									,.R1(R[491])	,.R2(R[634])									,.clk(clk)	,.L(L386)	,.P(P[385])	,.reset(reset)	);
VNU_2 VNU387	(.Q1(Q[497])	,.Q2(Q[640])									,.R1(R[497])	,.R2(R[640])									,.clk(clk)	,.L(L387)	,.P(P[386])	,.reset(reset)	);
VNU_2 VNU388	(.Q1(Q[503])	,.Q2(Q[646])									,.R1(R[503])	,.R2(R[646])									,.clk(clk)	,.L(L388)	,.P(P[387])	,.reset(reset)	);
VNU_2 VNU389	(.Q1(Q[509])	,.Q2(Q[652])									,.R1(R[509])	,.R2(R[652])									,.clk(clk)	,.L(L389)	,.P(P[388])	,.reset(reset)	);
VNU_2 VNU390	(.Q1(Q[515])	,.Q2(Q[658])									,.R1(R[515])	,.R2(R[658])									,.clk(clk)	,.L(L390)	,.P(P[389])	,.reset(reset)	);
VNU_2 VNU391	(.Q1(Q[521])	,.Q2(Q[664])									,.R1(R[521])	,.R2(R[664])									,.clk(clk)	,.L(L391)	,.P(P[390])	,.reset(reset)	);
VNU_2 VNU392	(.Q1(Q[527])	,.Q2(Q[670])									,.R1(R[527])	,.R2(R[670])									,.clk(clk)	,.L(L392)	,.P(P[391])	,.reset(reset)	);
VNU_2 VNU393	(.Q1(Q[533])	,.Q2(Q[676])									,.R1(R[533])	,.R2(R[676])									,.clk(clk)	,.L(L393)	,.P(P[392])	,.reset(reset)	);
VNU_2 VNU394	(.Q1(Q[539])	,.Q2(Q[682])									,.R1(R[539])	,.R2(R[682])									,.clk(clk)	,.L(L394)	,.P(P[393])	,.reset(reset)	);
VNU_2 VNU395	(.Q1(Q[545])	,.Q2(Q[688])									,.R1(R[545])	,.R2(R[688])									,.clk(clk)	,.L(L395)	,.P(P[394])	,.reset(reset)	);
VNU_2 VNU396	(.Q1(Q[551])	,.Q2(Q[694])									,.R1(R[551])	,.R2(R[694])									,.clk(clk)	,.L(L396)	,.P(P[395])	,.reset(reset)	);
VNU_2 VNU397	(.Q1(Q[557])	,.Q2(Q[700])									,.R1(R[557])	,.R2(R[700])									,.clk(clk)	,.L(L397)	,.P(P[396])	,.reset(reset)	);
VNU_2 VNU398	(.Q1(Q[563])	,.Q2(Q[706])									,.R1(R[563])	,.R2(R[706])									,.clk(clk)	,.L(L398)	,.P(P[397])	,.reset(reset)	);
VNU_2 VNU399	(.Q1(Q[569])	,.Q2(Q[712])									,.R1(R[569])	,.R2(R[712])									,.clk(clk)	,.L(L399)	,.P(P[398])	,.reset(reset)	);
VNU_2 VNU400	(.Q1(Q[575])	,.Q2(Q[718])									,.R1(R[575])	,.R2(R[718])									,.clk(clk)	,.L(L400)	,.P(P[399])	,.reset(reset)	);
VNU_2 VNU401	(.Q1(Q[581])	,.Q2(Q[724])									,.R1(R[581])	,.R2(R[724])									,.clk(clk)	,.L(L401)	,.P(P[400])	,.reset(reset)	);
VNU_2 VNU402	(.Q1(Q[587])	,.Q2(Q[730])									,.R1(R[587])	,.R2(R[730])									,.clk(clk)	,.L(L402)	,.P(P[401])	,.reset(reset)	);
VNU_2 VNU403	(.Q1(Q[593])	,.Q2(Q[736])									,.R1(R[593])	,.R2(R[736])									,.clk(clk)	,.L(L403)	,.P(P[402])	,.reset(reset)	);
VNU_2 VNU404	(.Q1(Q[599])	,.Q2(Q[742])									,.R1(R[599])	,.R2(R[742])									,.clk(clk)	,.L(L404)	,.P(P[403])	,.reset(reset)	);
VNU_2 VNU405	(.Q1(Q[605])	,.Q2(Q[748])									,.R1(R[605])	,.R2(R[748])									,.clk(clk)	,.L(L405)	,.P(P[404])	,.reset(reset)	);
VNU_2 VNU406	(.Q1(Q[611])	,.Q2(Q[754])									,.R1(R[611])	,.R2(R[754])									,.clk(clk)	,.L(L406)	,.P(P[405])	,.reset(reset)	);
VNU_2 VNU407	(.Q1(Q[617])	,.Q2(Q[760])									,.R1(R[617])	,.R2(R[760])									,.clk(clk)	,.L(L407)	,.P(P[406])	,.reset(reset)	);
VNU_2 VNU408	(.Q1(Q[623])	,.Q2(Q[766])									,.R1(R[623])	,.R2(R[766])									,.clk(clk)	,.L(L408)	,.P(P[407])	,.reset(reset)	);
VNU_2 VNU409	(.Q1(Q[629])	,.Q2(Q[773])									,.R1(R[629])	,.R2(R[773])									,.clk(clk)	,.L(L409)	,.P(P[408])	,.reset(reset)	);
VNU_2 VNU410	(.Q1(Q[635])	,.Q2(Q[780])									,.R1(R[635])	,.R2(R[780])									,.clk(clk)	,.L(L410)	,.P(P[409])	,.reset(reset)	);
VNU_2 VNU411	(.Q1(Q[641])	,.Q2(Q[787])									,.R1(R[641])	,.R2(R[787])									,.clk(clk)	,.L(L411)	,.P(P[410])	,.reset(reset)	);
VNU_2 VNU412	(.Q1(Q[647])	,.Q2(Q[794])									,.R1(R[647])	,.R2(R[794])									,.clk(clk)	,.L(L412)	,.P(P[411])	,.reset(reset)	);
VNU_2 VNU413	(.Q1(Q[653])	,.Q2(Q[801])									,.R1(R[653])	,.R2(R[801])									,.clk(clk)	,.L(L413)	,.P(P[412])	,.reset(reset)	);
VNU_2 VNU414	(.Q1(Q[659])	,.Q2(Q[808])									,.R1(R[659])	,.R2(R[808])									,.clk(clk)	,.L(L414)	,.P(P[413])	,.reset(reset)	);
VNU_2 VNU415	(.Q1(Q[665])	,.Q2(Q[815])									,.R1(R[665])	,.R2(R[815])									,.clk(clk)	,.L(L415)	,.P(P[414])	,.reset(reset)	);
VNU_2 VNU416	(.Q1(Q[671])	,.Q2(Q[822])									,.R1(R[671])	,.R2(R[822])									,.clk(clk)	,.L(L416)	,.P(P[415])	,.reset(reset)	);
VNU_2 VNU417	(.Q1(Q[677])	,.Q2(Q[829])									,.R1(R[677])	,.R2(R[829])									,.clk(clk)	,.L(L417)	,.P(P[416])	,.reset(reset)	);
VNU_2 VNU418	(.Q1(Q[683])	,.Q2(Q[836])									,.R1(R[683])	,.R2(R[836])									,.clk(clk)	,.L(L418)	,.P(P[417])	,.reset(reset)	);
VNU_2 VNU419	(.Q1(Q[689])	,.Q2(Q[843])									,.R1(R[689])	,.R2(R[843])									,.clk(clk)	,.L(L419)	,.P(P[418])	,.reset(reset)	);
VNU_2 VNU420	(.Q1(Q[695])	,.Q2(Q[850])									,.R1(R[695])	,.R2(R[850])									,.clk(clk)	,.L(L420)	,.P(P[419])	,.reset(reset)	);
VNU_2 VNU421	(.Q1(Q[701])	,.Q2(Q[857])									,.R1(R[701])	,.R2(R[857])									,.clk(clk)	,.L(L421)	,.P(P[420])	,.reset(reset)	);
VNU_2 VNU422	(.Q1(Q[707])	,.Q2(Q[864])									,.R1(R[707])	,.R2(R[864])									,.clk(clk)	,.L(L422)	,.P(P[421])	,.reset(reset)	);
VNU_2 VNU423	(.Q1(Q[713])	,.Q2(Q[871])									,.R1(R[713])	,.R2(R[871])									,.clk(clk)	,.L(L423)	,.P(P[422])	,.reset(reset)	);
VNU_2 VNU424	(.Q1(Q[719])	,.Q2(Q[878])									,.R1(R[719])	,.R2(R[878])									,.clk(clk)	,.L(L424)	,.P(P[423])	,.reset(reset)	);
VNU_2 VNU425	(.Q1(Q[725])	,.Q2(Q[885])									,.R1(R[725])	,.R2(R[885])									,.clk(clk)	,.L(L425)	,.P(P[424])	,.reset(reset)	);
VNU_2 VNU426	(.Q1(Q[731])	,.Q2(Q[892])									,.R1(R[731])	,.R2(R[892])									,.clk(clk)	,.L(L426)	,.P(P[425])	,.reset(reset)	);
VNU_2 VNU427	(.Q1(Q[737])	,.Q2(Q[899])									,.R1(R[737])	,.R2(R[899])									,.clk(clk)	,.L(L427)	,.P(P[426])	,.reset(reset)	);
VNU_2 VNU428	(.Q1(Q[743])	,.Q2(Q[906])									,.R1(R[743])	,.R2(R[906])									,.clk(clk)	,.L(L428)	,.P(P[427])	,.reset(reset)	);
VNU_2 VNU429	(.Q1(Q[749])	,.Q2(Q[913])									,.R1(R[749])	,.R2(R[913])									,.clk(clk)	,.L(L429)	,.P(P[428])	,.reset(reset)	);
VNU_2 VNU430	(.Q1(Q[755])	,.Q2(Q[920])									,.R1(R[755])	,.R2(R[920])									,.clk(clk)	,.L(L430)	,.P(P[429])	,.reset(reset)	);
VNU_2 VNU431	(.Q1(Q[761])	,.Q2(Q[927])									,.R1(R[761])	,.R2(R[927])									,.clk(clk)	,.L(L431)	,.P(P[430])	,.reset(reset)	);
VNU_2 VNU432	(.Q1(Q[767])	,.Q2(Q[934])									,.R1(R[767])	,.R2(R[934])									,.clk(clk)	,.L(L432)	,.P(P[431])	,.reset(reset)	);
VNU_2 VNU433	(.Q1(Q[774])	,.Q2(Q[940])									,.R1(R[774])	,.R2(R[940])									,.clk(clk)	,.L(L433)	,.P(P[432])	,.reset(reset)	);
VNU_2 VNU434	(.Q1(Q[781])	,.Q2(Q[946])									,.R1(R[781])	,.R2(R[946])									,.clk(clk)	,.L(L434)	,.P(P[433])	,.reset(reset)	);
VNU_2 VNU435	(.Q1(Q[788])	,.Q2(Q[952])									,.R1(R[788])	,.R2(R[952])									,.clk(clk)	,.L(L435)	,.P(P[434])	,.reset(reset)	);
VNU_2 VNU436	(.Q1(Q[795])	,.Q2(Q[958])									,.R1(R[795])	,.R2(R[958])									,.clk(clk)	,.L(L436)	,.P(P[435])	,.reset(reset)	);
VNU_2 VNU437	(.Q1(Q[802])	,.Q2(Q[964])									,.R1(R[802])	,.R2(R[964])									,.clk(clk)	,.L(L437)	,.P(P[436])	,.reset(reset)	);
VNU_2 VNU438	(.Q1(Q[809])	,.Q2(Q[970])									,.R1(R[809])	,.R2(R[970])									,.clk(clk)	,.L(L438)	,.P(P[437])	,.reset(reset)	);
VNU_2 VNU439	(.Q1(Q[816])	,.Q2(Q[976])									,.R1(R[816])	,.R2(R[976])									,.clk(clk)	,.L(L439)	,.P(P[438])	,.reset(reset)	);
VNU_2 VNU440	(.Q1(Q[823])	,.Q2(Q[982])									,.R1(R[823])	,.R2(R[982])									,.clk(clk)	,.L(L440)	,.P(P[439])	,.reset(reset)	);
VNU_2 VNU441	(.Q1(Q[830])	,.Q2(Q[988])									,.R1(R[830])	,.R2(R[988])									,.clk(clk)	,.L(L441)	,.P(P[440])	,.reset(reset)	);
VNU_2 VNU442	(.Q1(Q[837])	,.Q2(Q[994])									,.R1(R[837])	,.R2(R[994])									,.clk(clk)	,.L(L442)	,.P(P[441])	,.reset(reset)	);
VNU_2 VNU443	(.Q1(Q[844])	,.Q2(Q[1000])									,.R1(R[844])	,.R2(R[1000])									,.clk(clk)	,.L(L443)	,.P(P[442])	,.reset(reset)	);
VNU_2 VNU444	(.Q1(Q[851])	,.Q2(Q[1006])									,.R1(R[851])	,.R2(R[1006])									,.clk(clk)	,.L(L444)	,.P(P[443])	,.reset(reset)	);
VNU_2 VNU445	(.Q1(Q[858])	,.Q2(Q[1012])									,.R1(R[858])	,.R2(R[1012])									,.clk(clk)	,.L(L445)	,.P(P[444])	,.reset(reset)	);
VNU_2 VNU446	(.Q1(Q[865])	,.Q2(Q[1018])									,.R1(R[865])	,.R2(R[1018])									,.clk(clk)	,.L(L446)	,.P(P[445])	,.reset(reset)	);
VNU_2 VNU447	(.Q1(Q[872])	,.Q2(Q[1024])									,.R1(R[872])	,.R2(R[1024])									,.clk(clk)	,.L(L447)	,.P(P[446])	,.reset(reset)	);
VNU_2 VNU448	(.Q1(Q[879])	,.Q2(Q[1030])									,.R1(R[879])	,.R2(R[1030])									,.clk(clk)	,.L(L448)	,.P(P[447])	,.reset(reset)	);
VNU_2 VNU449	(.Q1(Q[886])	,.Q2(Q[1036])									,.R1(R[886])	,.R2(R[1036])									,.clk(clk)	,.L(L449)	,.P(P[448])	,.reset(reset)	);
VNU_2 VNU450	(.Q1(Q[893])	,.Q2(Q[1042])									,.R1(R[893])	,.R2(R[1042])									,.clk(clk)	,.L(L450)	,.P(P[449])	,.reset(reset)	);
VNU_2 VNU451	(.Q1(Q[900])	,.Q2(Q[1048])									,.R1(R[900])	,.R2(R[1048])									,.clk(clk)	,.L(L451)	,.P(P[450])	,.reset(reset)	);
VNU_2 VNU452	(.Q1(Q[907])	,.Q2(Q[1054])									,.R1(R[907])	,.R2(R[1054])									,.clk(clk)	,.L(L452)	,.P(P[451])	,.reset(reset)	);
VNU_2 VNU453	(.Q1(Q[914])	,.Q2(Q[1060])									,.R1(R[914])	,.R2(R[1060])									,.clk(clk)	,.L(L453)	,.P(P[452])	,.reset(reset)	);
VNU_2 VNU454	(.Q1(Q[921])	,.Q2(Q[1066])									,.R1(R[921])	,.R2(R[1066])									,.clk(clk)	,.L(L454)	,.P(P[453])	,.reset(reset)	);
VNU_2 VNU455	(.Q1(Q[928])	,.Q2(Q[1072])									,.R1(R[928])	,.R2(R[1072])									,.clk(clk)	,.L(L455)	,.P(P[454])	,.reset(reset)	);
VNU_2 VNU456	(.Q1(Q[935])	,.Q2(Q[1078])									,.R1(R[935])	,.R2(R[1078])									,.clk(clk)	,.L(L456)	,.P(P[455])	,.reset(reset)	);
VNU_2 VNU457	(.Q1(Q[941])	,.Q2(Q[1084])									,.R1(R[941])	,.R2(R[1084])									,.clk(clk)	,.L(L457)	,.P(P[456])	,.reset(reset)	);
VNU_2 VNU458	(.Q1(Q[947])	,.Q2(Q[1090])									,.R1(R[947])	,.R2(R[1090])									,.clk(clk)	,.L(L458)	,.P(P[457])	,.reset(reset)	);
VNU_2 VNU459	(.Q1(Q[953])	,.Q2(Q[1096])									,.R1(R[953])	,.R2(R[1096])									,.clk(clk)	,.L(L459)	,.P(P[458])	,.reset(reset)	);
VNU_2 VNU460	(.Q1(Q[959])	,.Q2(Q[1102])									,.R1(R[959])	,.R2(R[1102])									,.clk(clk)	,.L(L460)	,.P(P[459])	,.reset(reset)	);
VNU_2 VNU461	(.Q1(Q[965])	,.Q2(Q[1108])									,.R1(R[965])	,.R2(R[1108])									,.clk(clk)	,.L(L461)	,.P(P[460])	,.reset(reset)	);
VNU_2 VNU462	(.Q1(Q[971])	,.Q2(Q[1114])									,.R1(R[971])	,.R2(R[1114])									,.clk(clk)	,.L(L462)	,.P(P[461])	,.reset(reset)	);
VNU_2 VNU463	(.Q1(Q[977])	,.Q2(Q[1120])									,.R1(R[977])	,.R2(R[1120])									,.clk(clk)	,.L(L463)	,.P(P[462])	,.reset(reset)	);
VNU_2 VNU464	(.Q1(Q[983])	,.Q2(Q[1126])									,.R1(R[983])	,.R2(R[1126])									,.clk(clk)	,.L(L464)	,.P(P[463])	,.reset(reset)	);
VNU_2 VNU465	(.Q1(Q[989])	,.Q2(Q[1132])									,.R1(R[989])	,.R2(R[1132])									,.clk(clk)	,.L(L465)	,.P(P[464])	,.reset(reset)	);
VNU_2 VNU466	(.Q1(Q[995])	,.Q2(Q[1138])									,.R1(R[995])	,.R2(R[1138])									,.clk(clk)	,.L(L466)	,.P(P[465])	,.reset(reset)	);
VNU_2 VNU467	(.Q1(Q[1001])	,.Q2(Q[1144])									,.R1(R[1001])	,.R2(R[1144])									,.clk(clk)	,.L(L467)	,.P(P[466])	,.reset(reset)	);
VNU_2 VNU468	(.Q1(Q[1007])	,.Q2(Q[1150])									,.R1(R[1007])	,.R2(R[1150])									,.clk(clk)	,.L(L468)	,.P(P[467])	,.reset(reset)	);
VNU_2 VNU469	(.Q1(Q[1013])	,.Q2(Q[1156])									,.R1(R[1013])	,.R2(R[1156])									,.clk(clk)	,.L(L469)	,.P(P[468])	,.reset(reset)	);
VNU_2 VNU470	(.Q1(Q[1019])	,.Q2(Q[1162])									,.R1(R[1019])	,.R2(R[1162])									,.clk(clk)	,.L(L470)	,.P(P[469])	,.reset(reset)	);
VNU_2 VNU471	(.Q1(Q[1025])	,.Q2(Q[1168])									,.R1(R[1025])	,.R2(R[1168])									,.clk(clk)	,.L(L471)	,.P(P[470])	,.reset(reset)	);
VNU_2 VNU472	(.Q1(Q[1031])	,.Q2(Q[1174])									,.R1(R[1031])	,.R2(R[1174])									,.clk(clk)	,.L(L472)	,.P(P[471])	,.reset(reset)	);
VNU_2 VNU473	(.Q1(Q[1037])	,.Q2(Q[1180])									,.R1(R[1037])	,.R2(R[1180])									,.clk(clk)	,.L(L473)	,.P(P[472])	,.reset(reset)	);
VNU_2 VNU474	(.Q1(Q[1043])	,.Q2(Q[1186])									,.R1(R[1043])	,.R2(R[1186])									,.clk(clk)	,.L(L474)	,.P(P[473])	,.reset(reset)	);
VNU_2 VNU475	(.Q1(Q[1049])	,.Q2(Q[1192])									,.R1(R[1049])	,.R2(R[1192])									,.clk(clk)	,.L(L475)	,.P(P[474])	,.reset(reset)	);
VNU_2 VNU476	(.Q1(Q[1055])	,.Q2(Q[1198])									,.R1(R[1055])	,.R2(R[1198])									,.clk(clk)	,.L(L476)	,.P(P[475])	,.reset(reset)	);
VNU_2 VNU477	(.Q1(Q[1061])	,.Q2(Q[1204])									,.R1(R[1061])	,.R2(R[1204])									,.clk(clk)	,.L(L477)	,.P(P[476])	,.reset(reset)	);
VNU_2 VNU478	(.Q1(Q[1067])	,.Q2(Q[1210])									,.R1(R[1067])	,.R2(R[1210])									,.clk(clk)	,.L(L478)	,.P(P[477])	,.reset(reset)	);
VNU_2 VNU479	(.Q1(Q[1073])	,.Q2(Q[1216])									,.R1(R[1073])	,.R2(R[1216])									,.clk(clk)	,.L(L479)	,.P(P[478])	,.reset(reset)	);
VNU_2 VNU480	(.Q1(Q[1079])	,.Q2(Q[1222])									,.R1(R[1079])	,.R2(R[1222])									,.clk(clk)	,.L(L480)	,.P(P[479])	,.reset(reset)	);
VNU_2 VNU481	(.Q1(Q[1085])	,.Q2(Q[1229])									,.R1(R[1085])	,.R2(R[1229])									,.clk(clk)	,.L(L481)	,.P(P[480])	,.reset(reset)	);
VNU_2 VNU482	(.Q1(Q[1091])	,.Q2(Q[1236])									,.R1(R[1091])	,.R2(R[1236])									,.clk(clk)	,.L(L482)	,.P(P[481])	,.reset(reset)	);
VNU_2 VNU483	(.Q1(Q[1097])	,.Q2(Q[1243])									,.R1(R[1097])	,.R2(R[1243])									,.clk(clk)	,.L(L483)	,.P(P[482])	,.reset(reset)	);
VNU_2 VNU484	(.Q1(Q[1103])	,.Q2(Q[1250])									,.R1(R[1103])	,.R2(R[1250])									,.clk(clk)	,.L(L484)	,.P(P[483])	,.reset(reset)	);
VNU_2 VNU485	(.Q1(Q[1109])	,.Q2(Q[1257])									,.R1(R[1109])	,.R2(R[1257])									,.clk(clk)	,.L(L485)	,.P(P[484])	,.reset(reset)	);
VNU_2 VNU486	(.Q1(Q[1115])	,.Q2(Q[1264])									,.R1(R[1115])	,.R2(R[1264])									,.clk(clk)	,.L(L486)	,.P(P[485])	,.reset(reset)	);
VNU_2 VNU487	(.Q1(Q[1121])	,.Q2(Q[1271])									,.R1(R[1121])	,.R2(R[1271])									,.clk(clk)	,.L(L487)	,.P(P[486])	,.reset(reset)	);
VNU_2 VNU488	(.Q1(Q[1127])	,.Q2(Q[1278])									,.R1(R[1127])	,.R2(R[1278])									,.clk(clk)	,.L(L488)	,.P(P[487])	,.reset(reset)	);
VNU_2 VNU489	(.Q1(Q[1133])	,.Q2(Q[1285])									,.R1(R[1133])	,.R2(R[1285])									,.clk(clk)	,.L(L489)	,.P(P[488])	,.reset(reset)	);
VNU_2 VNU490	(.Q1(Q[1139])	,.Q2(Q[1292])									,.R1(R[1139])	,.R2(R[1292])									,.clk(clk)	,.L(L490)	,.P(P[489])	,.reset(reset)	);
VNU_2 VNU491	(.Q1(Q[1145])	,.Q2(Q[1299])									,.R1(R[1145])	,.R2(R[1299])									,.clk(clk)	,.L(L491)	,.P(P[490])	,.reset(reset)	);
VNU_2 VNU492	(.Q1(Q[1151])	,.Q2(Q[1306])									,.R1(R[1151])	,.R2(R[1306])									,.clk(clk)	,.L(L492)	,.P(P[491])	,.reset(reset)	);
VNU_2 VNU493	(.Q1(Q[1157])	,.Q2(Q[1313])									,.R1(R[1157])	,.R2(R[1313])									,.clk(clk)	,.L(L493)	,.P(P[492])	,.reset(reset)	);
VNU_2 VNU494	(.Q1(Q[1163])	,.Q2(Q[1320])									,.R1(R[1163])	,.R2(R[1320])									,.clk(clk)	,.L(L494)	,.P(P[493])	,.reset(reset)	);
VNU_2 VNU495	(.Q1(Q[1169])	,.Q2(Q[1327])									,.R1(R[1169])	,.R2(R[1327])									,.clk(clk)	,.L(L495)	,.P(P[494])	,.reset(reset)	);
VNU_2 VNU496	(.Q1(Q[1175])	,.Q2(Q[1334])									,.R1(R[1175])	,.R2(R[1334])									,.clk(clk)	,.L(L496)	,.P(P[495])	,.reset(reset)	);
VNU_2 VNU497	(.Q1(Q[1181])	,.Q2(Q[1341])									,.R1(R[1181])	,.R2(R[1341])									,.clk(clk)	,.L(L497)	,.P(P[496])	,.reset(reset)	);
VNU_2 VNU498	(.Q1(Q[1187])	,.Q2(Q[1348])									,.R1(R[1187])	,.R2(R[1348])									,.clk(clk)	,.L(L498)	,.P(P[497])	,.reset(reset)	);
VNU_2 VNU499	(.Q1(Q[1193])	,.Q2(Q[1355])									,.R1(R[1193])	,.R2(R[1355])									,.clk(clk)	,.L(L499)	,.P(P[498])	,.reset(reset)	);
VNU_2 VNU500	(.Q1(Q[1199])	,.Q2(Q[1362])									,.R1(R[1199])	,.R2(R[1362])									,.clk(clk)	,.L(L500)	,.P(P[499])	,.reset(reset)	);
VNU_2 VNU501	(.Q1(Q[1205])	,.Q2(Q[1369])									,.R1(R[1205])	,.R2(R[1369])									,.clk(clk)	,.L(L501)	,.P(P[500])	,.reset(reset)	);
VNU_2 VNU502	(.Q1(Q[1211])	,.Q2(Q[1376])									,.R1(R[1211])	,.R2(R[1376])									,.clk(clk)	,.L(L502)	,.P(P[501])	,.reset(reset)	);
VNU_2 VNU503	(.Q1(Q[1217])	,.Q2(Q[1383])									,.R1(R[1217])	,.R2(R[1383])									,.clk(clk)	,.L(L503)	,.P(P[502])	,.reset(reset)	);
VNU_2 VNU504	(.Q1(Q[1223])	,.Q2(Q[1390])									,.R1(R[1223])	,.R2(R[1390])									,.clk(clk)	,.L(L504)	,.P(P[503])	,.reset(reset)	);
VNU_2 VNU505	(.Q1(Q[1230])	,.Q2(Q[1396])									,.R1(R[1230])	,.R2(R[1396])									,.clk(clk)	,.L(L505)	,.P(P[504])	,.reset(reset)	);
VNU_2 VNU506	(.Q1(Q[1237])	,.Q2(Q[1402])									,.R1(R[1237])	,.R2(R[1402])									,.clk(clk)	,.L(L506)	,.P(P[505])	,.reset(reset)	);
VNU_2 VNU507	(.Q1(Q[1244])	,.Q2(Q[1408])									,.R1(R[1244])	,.R2(R[1408])									,.clk(clk)	,.L(L507)	,.P(P[506])	,.reset(reset)	);
VNU_2 VNU508	(.Q1(Q[1251])	,.Q2(Q[1414])									,.R1(R[1251])	,.R2(R[1414])									,.clk(clk)	,.L(L508)	,.P(P[507])	,.reset(reset)	);
VNU_2 VNU509	(.Q1(Q[1258])	,.Q2(Q[1420])									,.R1(R[1258])	,.R2(R[1420])									,.clk(clk)	,.L(L509)	,.P(P[508])	,.reset(reset)	);
VNU_2 VNU510	(.Q1(Q[1265])	,.Q2(Q[1426])									,.R1(R[1265])	,.R2(R[1426])									,.clk(clk)	,.L(L510)	,.P(P[509])	,.reset(reset)	);
VNU_2 VNU511	(.Q1(Q[1272])	,.Q2(Q[1432])									,.R1(R[1272])	,.R2(R[1432])									,.clk(clk)	,.L(L511)	,.P(P[510])	,.reset(reset)	);
VNU_2 VNU512	(.Q1(Q[1279])	,.Q2(Q[1438])									,.R1(R[1279])	,.R2(R[1438])									,.clk(clk)	,.L(L512)	,.P(P[511])	,.reset(reset)	);
VNU_2 VNU513	(.Q1(Q[1286])	,.Q2(Q[1444])									,.R1(R[1286])	,.R2(R[1444])									,.clk(clk)	,.L(L513)	,.P(P[512])	,.reset(reset)	);
VNU_2 VNU514	(.Q1(Q[1293])	,.Q2(Q[1450])									,.R1(R[1293])	,.R2(R[1450])									,.clk(clk)	,.L(L514)	,.P(P[513])	,.reset(reset)	);
VNU_2 VNU515	(.Q1(Q[1300])	,.Q2(Q[1456])									,.R1(R[1300])	,.R2(R[1456])									,.clk(clk)	,.L(L515)	,.P(P[514])	,.reset(reset)	);
VNU_2 VNU516	(.Q1(Q[1307])	,.Q2(Q[1462])									,.R1(R[1307])	,.R2(R[1462])									,.clk(clk)	,.L(L516)	,.P(P[515])	,.reset(reset)	);
VNU_2 VNU517	(.Q1(Q[1314])	,.Q2(Q[1468])									,.R1(R[1314])	,.R2(R[1468])									,.clk(clk)	,.L(L517)	,.P(P[516])	,.reset(reset)	);
VNU_2 VNU518	(.Q1(Q[1321])	,.Q2(Q[1474])									,.R1(R[1321])	,.R2(R[1474])									,.clk(clk)	,.L(L518)	,.P(P[517])	,.reset(reset)	);
VNU_2 VNU519	(.Q1(Q[1328])	,.Q2(Q[1480])									,.R1(R[1328])	,.R2(R[1480])									,.clk(clk)	,.L(L519)	,.P(P[518])	,.reset(reset)	);
VNU_2 VNU520	(.Q1(Q[1335])	,.Q2(Q[1486])									,.R1(R[1335])	,.R2(R[1486])									,.clk(clk)	,.L(L520)	,.P(P[519])	,.reset(reset)	);
VNU_2 VNU521	(.Q1(Q[1342])	,.Q2(Q[1492])									,.R1(R[1342])	,.R2(R[1492])									,.clk(clk)	,.L(L521)	,.P(P[520])	,.reset(reset)	);
VNU_2 VNU522	(.Q1(Q[1349])	,.Q2(Q[1498])									,.R1(R[1349])	,.R2(R[1498])									,.clk(clk)	,.L(L522)	,.P(P[521])	,.reset(reset)	);
VNU_2 VNU523	(.Q1(Q[1356])	,.Q2(Q[1504])									,.R1(R[1356])	,.R2(R[1504])									,.clk(clk)	,.L(L523)	,.P(P[522])	,.reset(reset)	);
VNU_2 VNU524	(.Q1(Q[1363])	,.Q2(Q[1510])									,.R1(R[1363])	,.R2(R[1510])									,.clk(clk)	,.L(L524)	,.P(P[523])	,.reset(reset)	);
VNU_2 VNU525	(.Q1(Q[1370])	,.Q2(Q[1516])									,.R1(R[1370])	,.R2(R[1516])									,.clk(clk)	,.L(L525)	,.P(P[524])	,.reset(reset)	);
VNU_2 VNU526	(.Q1(Q[1377])	,.Q2(Q[1522])									,.R1(R[1377])	,.R2(R[1522])									,.clk(clk)	,.L(L526)	,.P(P[525])	,.reset(reset)	);
VNU_2 VNU527	(.Q1(Q[1384])	,.Q2(Q[1528])									,.R1(R[1384])	,.R2(R[1528])									,.clk(clk)	,.L(L527)	,.P(P[526])	,.reset(reset)	);
VNU_2 VNU528	(.Q1(Q[1391])	,.Q2(Q[1534])									,.R1(R[1391])	,.R2(R[1534])									,.clk(clk)	,.L(L528)	,.P(P[527])	,.reset(reset)	);
VNU_2 VNU529	(.Q1(Q[1397])	,.Q2(Q[1540])									,.R1(R[1397])	,.R2(R[1540])									,.clk(clk)	,.L(L529)	,.P(P[528])	,.reset(reset)	);
VNU_2 VNU530	(.Q1(Q[1403])	,.Q2(Q[1546])									,.R1(R[1403])	,.R2(R[1546])									,.clk(clk)	,.L(L530)	,.P(P[529])	,.reset(reset)	);
VNU_2 VNU531	(.Q1(Q[1409])	,.Q2(Q[1552])									,.R1(R[1409])	,.R2(R[1552])									,.clk(clk)	,.L(L531)	,.P(P[530])	,.reset(reset)	);
VNU_2 VNU532	(.Q1(Q[1415])	,.Q2(Q[1558])									,.R1(R[1415])	,.R2(R[1558])									,.clk(clk)	,.L(L532)	,.P(P[531])	,.reset(reset)	);
VNU_2 VNU533	(.Q1(Q[1421])	,.Q2(Q[1564])									,.R1(R[1421])	,.R2(R[1564])									,.clk(clk)	,.L(L533)	,.P(P[532])	,.reset(reset)	);
VNU_2 VNU534	(.Q1(Q[1427])	,.Q2(Q[1570])									,.R1(R[1427])	,.R2(R[1570])									,.clk(clk)	,.L(L534)	,.P(P[533])	,.reset(reset)	);
VNU_2 VNU535	(.Q1(Q[1433])	,.Q2(Q[1576])									,.R1(R[1433])	,.R2(R[1576])									,.clk(clk)	,.L(L535)	,.P(P[534])	,.reset(reset)	);
VNU_2 VNU536	(.Q1(Q[1439])	,.Q2(Q[1582])									,.R1(R[1439])	,.R2(R[1582])									,.clk(clk)	,.L(L536)	,.P(P[535])	,.reset(reset)	);
VNU_2 VNU537	(.Q1(Q[1445])	,.Q2(Q[1588])									,.R1(R[1445])	,.R2(R[1588])									,.clk(clk)	,.L(L537)	,.P(P[536])	,.reset(reset)	);
VNU_2 VNU538	(.Q1(Q[1451])	,.Q2(Q[1594])									,.R1(R[1451])	,.R2(R[1594])									,.clk(clk)	,.L(L538)	,.P(P[537])	,.reset(reset)	);
VNU_2 VNU539	(.Q1(Q[1457])	,.Q2(Q[1600])									,.R1(R[1457])	,.R2(R[1600])									,.clk(clk)	,.L(L539)	,.P(P[538])	,.reset(reset)	);
VNU_2 VNU540	(.Q1(Q[1463])	,.Q2(Q[1606])									,.R1(R[1463])	,.R2(R[1606])									,.clk(clk)	,.L(L540)	,.P(P[539])	,.reset(reset)	);
VNU_2 VNU541	(.Q1(Q[1469])	,.Q2(Q[1612])									,.R1(R[1469])	,.R2(R[1612])									,.clk(clk)	,.L(L541)	,.P(P[540])	,.reset(reset)	);
VNU_2 VNU542	(.Q1(Q[1475])	,.Q2(Q[1618])									,.R1(R[1475])	,.R2(R[1618])									,.clk(clk)	,.L(L542)	,.P(P[541])	,.reset(reset)	);
VNU_2 VNU543	(.Q1(Q[1481])	,.Q2(Q[1624])									,.R1(R[1481])	,.R2(R[1624])									,.clk(clk)	,.L(L543)	,.P(P[542])	,.reset(reset)	);
VNU_2 VNU544	(.Q1(Q[1487])	,.Q2(Q[1630])									,.R1(R[1487])	,.R2(R[1630])									,.clk(clk)	,.L(L544)	,.P(P[543])	,.reset(reset)	);
VNU_2 VNU545	(.Q1(Q[1493])	,.Q2(Q[1636])									,.R1(R[1493])	,.R2(R[1636])									,.clk(clk)	,.L(L545)	,.P(P[544])	,.reset(reset)	);
VNU_2 VNU546	(.Q1(Q[1499])	,.Q2(Q[1642])									,.R1(R[1499])	,.R2(R[1642])									,.clk(clk)	,.L(L546)	,.P(P[545])	,.reset(reset)	);
VNU_2 VNU547	(.Q1(Q[1505])	,.Q2(Q[1648])									,.R1(R[1505])	,.R2(R[1648])									,.clk(clk)	,.L(L547)	,.P(P[546])	,.reset(reset)	);
VNU_2 VNU548	(.Q1(Q[1511])	,.Q2(Q[1654])									,.R1(R[1511])	,.R2(R[1654])									,.clk(clk)	,.L(L548)	,.P(P[547])	,.reset(reset)	);
VNU_2 VNU549	(.Q1(Q[1517])	,.Q2(Q[1660])									,.R1(R[1517])	,.R2(R[1660])									,.clk(clk)	,.L(L549)	,.P(P[548])	,.reset(reset)	);
VNU_2 VNU550	(.Q1(Q[1523])	,.Q2(Q[1666])									,.R1(R[1523])	,.R2(R[1666])									,.clk(clk)	,.L(L550)	,.P(P[549])	,.reset(reset)	);
VNU_2 VNU551	(.Q1(Q[1529])	,.Q2(Q[1672])									,.R1(R[1529])	,.R2(R[1672])									,.clk(clk)	,.L(L551)	,.P(P[550])	,.reset(reset)	);
VNU_2 VNU552	(.Q1(Q[1535])	,.Q2(Q[1678])									,.R1(R[1535])	,.R2(R[1678])									,.clk(clk)	,.L(L552)	,.P(P[551])	,.reset(reset)	);
VNU_2 VNU553	(.Q1(Q[1541])	,.Q2(Q[1685])									,.R1(R[1541])	,.R2(R[1685])									,.clk(clk)	,.L(L553)	,.P(P[552])	,.reset(reset)	);
VNU_2 VNU554	(.Q1(Q[1547])	,.Q2(Q[1691])									,.R1(R[1547])	,.R2(R[1691])									,.clk(clk)	,.L(L554)	,.P(P[553])	,.reset(reset)	);
VNU_2 VNU555	(.Q1(Q[1553])	,.Q2(Q[1697])									,.R1(R[1553])	,.R2(R[1697])									,.clk(clk)	,.L(L555)	,.P(P[554])	,.reset(reset)	);
VNU_2 VNU556	(.Q1(Q[1559])	,.Q2(Q[1703])									,.R1(R[1559])	,.R2(R[1703])									,.clk(clk)	,.L(L556)	,.P(P[555])	,.reset(reset)	);
VNU_2 VNU557	(.Q1(Q[1565])	,.Q2(Q[1709])									,.R1(R[1565])	,.R2(R[1709])									,.clk(clk)	,.L(L557)	,.P(P[556])	,.reset(reset)	);
VNU_2 VNU558	(.Q1(Q[1571])	,.Q2(Q[1715])									,.R1(R[1571])	,.R2(R[1715])									,.clk(clk)	,.L(L558)	,.P(P[557])	,.reset(reset)	);
VNU_2 VNU559	(.Q1(Q[1577])	,.Q2(Q[1721])									,.R1(R[1577])	,.R2(R[1721])									,.clk(clk)	,.L(L559)	,.P(P[558])	,.reset(reset)	);
VNU_2 VNU560	(.Q1(Q[1583])	,.Q2(Q[1727])									,.R1(R[1583])	,.R2(R[1727])									,.clk(clk)	,.L(L560)	,.P(P[559])	,.reset(reset)	);
VNU_2 VNU561	(.Q1(Q[1589])	,.Q2(Q[1733])									,.R1(R[1589])	,.R2(R[1733])									,.clk(clk)	,.L(L561)	,.P(P[560])	,.reset(reset)	);
VNU_2 VNU562	(.Q1(Q[1595])	,.Q2(Q[1739])									,.R1(R[1595])	,.R2(R[1739])									,.clk(clk)	,.L(L562)	,.P(P[561])	,.reset(reset)	);
VNU_2 VNU563	(.Q1(Q[1601])	,.Q2(Q[1745])									,.R1(R[1601])	,.R2(R[1745])									,.clk(clk)	,.L(L563)	,.P(P[562])	,.reset(reset)	);
VNU_2 VNU564	(.Q1(Q[1607])	,.Q2(Q[1751])									,.R1(R[1607])	,.R2(R[1751])									,.clk(clk)	,.L(L564)	,.P(P[563])	,.reset(reset)	);
VNU_2 VNU565	(.Q1(Q[1613])	,.Q2(Q[1757])									,.R1(R[1613])	,.R2(R[1757])									,.clk(clk)	,.L(L565)	,.P(P[564])	,.reset(reset)	);
VNU_2 VNU566	(.Q1(Q[1619])	,.Q2(Q[1763])									,.R1(R[1619])	,.R2(R[1763])									,.clk(clk)	,.L(L566)	,.P(P[565])	,.reset(reset)	);
VNU_2 VNU567	(.Q1(Q[1625])	,.Q2(Q[1769])									,.R1(R[1625])	,.R2(R[1769])									,.clk(clk)	,.L(L567)	,.P(P[566])	,.reset(reset)	);
VNU_2 VNU568	(.Q1(Q[1631])	,.Q2(Q[1775])									,.R1(R[1631])	,.R2(R[1775])									,.clk(clk)	,.L(L568)	,.P(P[567])	,.reset(reset)	);
VNU_2 VNU569	(.Q1(Q[1637])	,.Q2(Q[1781])									,.R1(R[1637])	,.R2(R[1781])									,.clk(clk)	,.L(L569)	,.P(P[568])	,.reset(reset)	);
VNU_2 VNU570	(.Q1(Q[1643])	,.Q2(Q[1787])									,.R1(R[1643])	,.R2(R[1787])									,.clk(clk)	,.L(L570)	,.P(P[569])	,.reset(reset)	);
VNU_2 VNU571	(.Q1(Q[1649])	,.Q2(Q[1793])									,.R1(R[1649])	,.R2(R[1793])									,.clk(clk)	,.L(L571)	,.P(P[570])	,.reset(reset)	);
VNU_2 VNU572	(.Q1(Q[1655])	,.Q2(Q[1799])									,.R1(R[1655])	,.R2(R[1799])									,.clk(clk)	,.L(L572)	,.P(P[571])	,.reset(reset)	);
VNU_2 VNU573	(.Q1(Q[1661])	,.Q2(Q[1805])									,.R1(R[1661])	,.R2(R[1805])									,.clk(clk)	,.L(L573)	,.P(P[572])	,.reset(reset)	);
VNU_2 VNU574	(.Q1(Q[1667])	,.Q2(Q[1811])									,.R1(R[1667])	,.R2(R[1811])									,.clk(clk)	,.L(L574)	,.P(P[573])	,.reset(reset)	);
VNU_2 VNU575	(.Q1(Q[1673])	,.Q2(Q[1817])									,.R1(R[1673])	,.R2(R[1817])									,.clk(clk)	,.L(L575)	,.P(P[574])	,.reset(reset)	);
VNU_2 VNU576	(.Q1(Q[1679])	,.Q2(Q[1823])									,.R1(R[1679])	,.R2(R[1823])									,.clk(clk)	,.L(L576)	,.P(P[575])	,.reset(reset)	);

endmodule
